module sdoku_graph_mod (clk, rst, x, y, key, key_pulse,rgb,complete);


parameter X0 = 0;
parameter X1 = 71;
parameter X2 = 142;
parameter X3 = 213;
parameter X4 = 284;
parameter X5 = 355;
parameter X6 = 426;
parameter X7 = 497;
parameter X8 = 568;

parameter Y0 = 0;
parameter Y1 = 53;
parameter Y2 = 106;
parameter Y3 = 160;
parameter Y4 = 213;
parameter Y5 = 266;
parameter Y6 = 320;
parameter Y7 = 373;
parameter Y8 = 426;

input clk, rst;
input [9:0] x, y;
input [4:0] key, key_pulse; 
output [2:0]rgb;
output reg [1:0] complete;

wire [323:0] array;
wire line_on_h;
wire line_on_w;
wire line_on_bh;
wire line_on_bw;
wire [3:0] n;
wire [3:0] edit_x;
wire [3:0] edit_y;
wire [80:0] num;
wire [4:1] line1;
wire complete_tmp;


//module get_edit_n(input clk, rst, [4:0] key_pulse, 
//output reg [3:0] n, reg [3:0] edit_x,reg [3:0] edit_y);
get_edit_n d1(clk, rst, key_pulse,n,edit_x,edit_y);

//module number_input_mode1(input clk, rst , [4:0] key_pulse, [3:0] edit_x, [3:0] edit_y, [9:0]x, [9:0]y, [3:0] n,
// output reg[323:0] array);
number_input_mode1 d2(clk, rst, key_pulse, edit_x,edit_y,x,y,n,array);

//module complete_mode1(input clk, rst, [323:0] array , output check_tmp);
complete_mode1 d3 (clk, rst,key_pulse ,array,complete_tmp);


always@(*) begin
    case(complete_tmp)
       1'b0: complete = 2'b00;
       1'b1: complete = 2'b01;
       default : complete = 2'b11;
    endcase
end
                        
assign line_on_h = (x==71) || (x==142) ||  (x==284) || (x==355) || (x==497) || (x==568);
assign line_on_w = (y==53) || (y==106) || (y==213) || (y==266) || (y==373) || (y==426);

assign line_on_bh = (x >= 212 && x<= 214) || (x>=425 && x<= 427);
assign line_on_bw = (y>=159 && y<=161) || (y>=319 && y<=321);


 assign rgb =    cursor ? 3'b010 :
                (num[0]) ? 3'b001 :
                (num[1]) ? 3'b001 :
                (num[2]) ? 3'b000 :
                (num[3]) ? 3'b000 :
                (num[4]) ? 3'b001 :
                (num[5]) ? 3'b000 :
                (num[6]) ? 3'b000 :
                (num[7]) ? 3'b000 :
                (num[8]) ? 3'b000 :
                (num[9]) ? 3'b001 :
                (num[10]) ? 3'b000 :
                (num[11]) ? 3'b000 :
                (num[12]) ? 3'b001 :
                (num[13]) ? 3'b001 :
                (num[14]) ? 3'b001 :
                (num[15]) ? 3'b000 :
                (num[16]) ? 3'b000 :
                (num[17]) ? 3'b000 :
                (num[18]) ? 3'b000 :
                (num[19]) ? 3'b001 :
                (num[20]) ? 3'b001 :
                (num[21]) ? 3'b000 :
                (num[22]) ? 3'b000 :
                (num[23]) ? 3'b000 :
                (num[24]) ? 3'b000 :
                (num[25]) ? 3'b001 :
                (num[26]) ? 3'b000 :
                (num[27]) ? 3'b001 :
                (num[28]) ? 3'b000 :
                (num[29]) ? 3'b000 :
                (num[30]) ? 3'b000 :
                (num[31]) ? 3'b001 :
                (num[32]) ? 3'b000 :
                (num[33]) ? 3'b000 :
                (num[34]) ? 3'b000 :
                (num[35]) ? 3'b001 :
                (num[36]) ? 3'b001 :
                (num[37]) ? 3'b000 :
                (num[38]) ? 3'b000 :
                (num[39]) ? 3'b001 :
                (num[40]) ? 3'b000 :
                (num[41]) ? 3'b001 :
                (num[42]) ? 3'b000 :
                (num[43]) ? 3'b000 :
                (num[44]) ? 3'b001 :
                (num[45]) ? 3'b001 :
                (num[46]) ? 3'b000 :
                (num[47]) ? 3'b000 :
                (num[48]) ? 3'b000 :
                (num[49]) ? 3'b001 :
                (num[50]) ? 3'b000 :
                (num[51]) ? 3'b000 :
                (num[52]) ? 3'b000 :
                (num[53]) ? 3'b001 :
                (num[54]) ? 3'b000 :
                (num[55]) ? 3'b001 :
                (num[56]) ? 3'b000 :
                (num[57]) ? 3'b000 :
                (num[58]) ? 3'b000 :
                (num[59]) ? 3'b000 :
                (num[60]) ? 3'b001 :
                (num[61]) ? 3'b001 :
                (num[62]) ? 3'b000 :
                (num[63]) ? 3'b000 :
                (num[64]) ? 3'b000 :
                (num[65]) ? 3'b000 :
                (num[66]) ? 3'b001 :
                (num[67]) ? 3'b001 :
                (num[68]) ? 3'b001 :
                (num[69]) ? 3'b000 :
                (num[70]) ? 3'b000 :
                (num[71]) ? 3'b001 :
                (num[72]) ? 3'b000 :
                (num[73]) ? 3'b000 :
                (num[74]) ? 3'b000 :
                (num[75]) ? 3'b000 :
                (num[76]) ? 3'b001 :
                (num[77]) ? 3'b000 :
                (num[78]) ? 3'b000 :
                (num[79]) ? 3'b001 :
                (num[80]) ? 3'b001 :
                (line_on_bw) ? 3'b000 :
                (line_on_bh) ? 3'b000 : 
                (line_on_h) ? 3'b000 :
                (line_on_w) ? 3'b000 :
         
                3'b111;
               
 ///////////////////////////cursor//////////////////////////
  assign cursor = (edit_x == 0 && edit_y == 0) ? ((X0 + 11 < x && x < X0 + 56) && Y0 + 47 == y) :
                (edit_x == 1 && edit_y == 0) ? ((X1 + 11 < x && x < X1 + 56) && Y0 + 47 == y) :
                (edit_x == 2 && edit_y == 0) ? ((X2 + 11 < x && x < X2 + 56) && Y0 + 47 == y) :
                (edit_x == 3 && edit_y == 0) ? ((X3 + 11 < x && x < X3 + 56) && Y0 + 47 == y) :
                (edit_x == 4 && edit_y == 0) ? ((X4 + 11 < x && x < X4 + 56) && Y0 + 47 == y) :
                (edit_x == 5 && edit_y == 0) ? ((X5 + 11 < x && x < X5 + 56) && Y0 + 47 == y) :
                (edit_x == 6 && edit_y == 0) ? ((X6 + 11 < x && x < X6 + 56) && Y0 + 47 == y) :
                (edit_x == 7 && edit_y == 0) ? ((X7 + 11 < x && x < X7 + 56) && Y0 + 47 == y) :
                (edit_x == 8 && edit_y == 0) ? ((X8 + 11 < x && x < X8 + 56) && Y0 + 47 == y) :
                
                (edit_x == 0 && edit_y == 1) ? ((X0 + 11 < x && x < X0 + 56) && Y1 + 47 == y) :
                (edit_x == 1 && edit_y == 1) ? ((X1 + 11 < x && x < X1 + 56) && Y1 + 47 == y) :
                (edit_x == 2 && edit_y == 1) ? ((X2 + 11 < x && x < X2 + 56) && Y1 + 47 == y) :
                (edit_x == 3 && edit_y == 1) ? ((X3 + 11 < x && x < X3 + 56) && Y1 + 47 == y) :
                (edit_x == 4 && edit_y == 1) ? ((X4 + 11 < x && x < X4 + 56) && Y1 + 47 == y) :
                (edit_x == 5 && edit_y == 1) ? ((X5 + 11 < x && x < X5 + 56) && Y1 + 47 == y) :
                (edit_x == 6 && edit_y == 1) ? ((X6 + 11 < x && x < X6 + 56) && Y1 + 47 == y) :
                (edit_x == 7 && edit_y == 1) ? ((X7 + 11 < x && x < X7 + 56) && Y1 + 47 == y) :
                (edit_x == 8 && edit_y == 1) ? ((X8 + 11 < x && x < X8 + 56) && Y1 + 47 == y) :
                
                (edit_x == 0 && edit_y == 2) ? ((X0 + 11 < x && x < X0 + 56) && Y2 + 47 == y) :
                (edit_x == 1 && edit_y == 2) ? ((X1 + 11 < x && x < X1 + 56) && Y2 + 47 == y) :
                (edit_x == 2 && edit_y == 2) ? ((X2 + 11 < x && x < X2 + 56) && Y2 + 47 == y) :
                (edit_x == 3 && edit_y == 2) ? ((X3 + 11 < x && x < X3 + 56) && Y2 + 47 == y) :
                (edit_x == 4 && edit_y == 2) ? ((X4 + 11 < x && x < X4 + 56) && Y2 + 47 == y) :
                (edit_x == 5 && edit_y == 2) ? ((X5 + 11 < x && x < X5 + 56) && Y2 + 47 == y) :
                (edit_x == 6 && edit_y == 2) ? ((X6 + 11 < x && x < X6 + 56) && Y2 + 47 == y) :
                (edit_x == 7 && edit_y == 2) ? ((X7 + 11 < x && x < X7 + 56) && Y2 + 47 == y) :
                (edit_x == 8 && edit_y == 2) ? ((X8 + 11 < x && x < X8 + 56) && Y2 + 47 == y) :
                
                (edit_x == 0 && edit_y == 3) ? ((X0 + 11 < x && x < X0 + 56) && Y3 + 47 == y) :
                (edit_x == 1 && edit_y == 3) ? ((X1 + 11 < x && x < X1 + 56) && Y3 + 47 == y) :
                (edit_x == 2 && edit_y == 3) ? ((X2 + 11 < x && x < X2 + 56) && Y3 + 47 == y) :
                (edit_x == 3 && edit_y == 3) ? ((X3 + 11 < x && x < X3 + 56) && Y3 + 47 == y) :
                (edit_x == 4 && edit_y == 3) ? ((X4 + 11 < x && x < X4 + 56) && Y3 + 47 == y) :
                (edit_x == 5 && edit_y == 3) ? ((X5 + 11 < x && x < X5 + 56) && Y3 + 47 == y) :
                (edit_x == 6 && edit_y == 3) ? ((X6 + 11 < x && x < X6 + 56) && Y3 + 47 == y) :
                (edit_x == 7 && edit_y == 3) ? ((X7 + 11 < x && x < X7 + 56) && Y3 + 47 == y) :
                (edit_x == 8 && edit_y == 3) ? ((X8 + 11 < x && x < X8 + 56) && Y3 + 47 == y) :
                
                (edit_x == 0 && edit_y == 4) ? ((X0 + 11 < x && x < X0 + 56) && Y4 + 47 == y) :
                (edit_x == 1 && edit_y == 4) ? ((X1 + 11 < x && x < X1 + 56) && Y4 + 47 == y) :
                (edit_x == 2 && edit_y == 4) ? ((X2 + 11 < x && x < X2 + 56) && Y4 + 47 == y) :
                (edit_x == 3 && edit_y == 4) ? ((X3 + 11 < x && x < X3 + 56) && Y4 + 47 == y) :
                (edit_x == 4 && edit_y == 4) ? ((X4 + 11 < x && x < X4 + 56) && Y4 + 47 == y) :
                (edit_x == 5 && edit_y == 4) ? ((X5 + 11 < x && x < X5 + 56) && Y4 + 47 == y) :
                (edit_x == 6 && edit_y == 4) ? ((X6 + 11 < x && x < X6 + 56) && Y4 + 47 == y) :
                (edit_x == 7 && edit_y == 4) ? ((X7 + 11 < x && x < X7 + 56) && Y4 + 47 == y) :
                (edit_x == 8 && edit_y == 4) ? ((X8 + 11 < x && x < X8 + 56) && Y4 + 47 == y) :
                
                (edit_x == 0 && edit_y == 5) ? ((X0 + 11 < x && x < X0 + 56) && Y5 + 47 == y) :
                (edit_x == 1 && edit_y == 5) ? ((X1 + 11 < x && x < X1 + 56) && Y5 + 47 == y) :
                (edit_x == 2 && edit_y == 5) ? ((X2 + 11 < x && x < X2 + 56) && Y5 + 47 == y) :
                (edit_x == 3 && edit_y == 5) ? ((X3 + 11 < x && x < X3 + 56) && Y5 + 47 == y) :
                (edit_x == 4 && edit_y == 5) ? ((X4 + 11 < x && x < X4 + 56) && Y5 + 47 == y) :
                (edit_x == 5 && edit_y == 5) ? ((X5 + 11 < x && x < X5 + 56) && Y5 + 47 == y) :
                (edit_x == 6 && edit_y == 5) ? ((X6 + 11 < x && x < X6 + 56) && Y5 + 47 == y) :
                (edit_x == 7 && edit_y == 5) ? ((X7 + 11 < x && x < X7 + 56) && Y5 + 47 == y) :
                (edit_x == 8 && edit_y == 5) ? ((X8 + 11 < x && x < X8 + 56) && Y5 + 47 == y) :
                
                (edit_x == 0 && edit_y == 6) ? ((X0 + 11 < x && x < X0 + 56) && Y6 + 47 == y) :
                (edit_x == 1 && edit_y == 6) ? ((X1 + 11 < x && x < X1 + 56) && Y6 + 47 == y) :
                (edit_x == 2 && edit_y == 6) ? ((X2 + 11 < x && x < X2 + 56) && Y6 + 47 == y) :
                (edit_x == 3 && edit_y == 6) ? ((X3 + 11 < x && x < X3 + 56) && Y6 + 47 == y) :
                (edit_x == 4 && edit_y == 6) ? ((X4 + 11 < x && x < X4 + 56) && Y6 + 47 == y) :
                (edit_x == 5 && edit_y == 6) ? ((X5 + 11 < x && x < X5 + 56) && Y6 + 47 == y) :
                (edit_x == 6 && edit_y == 6) ? ((X6 + 11 < x && x < X6 + 56) && Y6 + 47 == y) :
                (edit_x == 7 && edit_y == 6) ? ((X7 + 11 < x && x < X7 + 56) && Y6 + 47 == y) :
                (edit_x == 8 && edit_y == 6) ? ((X8 + 11 < x && x < X8 + 56) && Y6 + 47 == y) :
                
                (edit_x == 0 && edit_y == 7) ? ((X0 + 11 < x && x < X0 + 56) && Y7 + 47 == y) :
                (edit_x == 1 && edit_y == 7) ? ((X1 + 11 < x && x < X1 + 56) && Y7 + 47 == y) :
                (edit_x == 2 && edit_y == 7) ? ((X2 + 11 < x && x < X2 + 56) && Y7 + 47 == y) :
                (edit_x == 3 && edit_y == 7) ? ((X3 + 11 < x && x < X3 + 56) && Y7 + 47 == y) :
                (edit_x == 4 && edit_y == 7) ? ((X4 + 11 < x && x < X4 + 56) && Y7 + 47 == y) :
                (edit_x == 5 && edit_y == 7) ? ((X5 + 11 < x && x < X5 + 56) && Y7 + 47 == y) :
                (edit_x == 6 && edit_y == 7) ? ((X6 + 11 < x && x < X6 + 56) && Y7 + 47 == y) :
                (edit_x == 7 && edit_y == 7) ? ((X7 + 11 < x && x < X7 + 56) && Y7 + 47 == y) :
                (edit_x == 8 && edit_y == 7) ? ((X8 + 11 < x && x < X8 + 56) && Y7 + 47 == y) :
                
                (edit_x == 0 && edit_y == 8) ? ((X0 + 11 < x && x < X0 + 56) && Y8 + 47 == y) :
                (edit_x == 1 && edit_y == 8) ? ((X1 + 11 < x && x < X1 + 56) && Y8 + 47 == y) :
                (edit_x == 2 && edit_y == 8) ? ((X2 + 11 < x && x < X2 + 56) && Y8 + 47 == y) :
                (edit_x == 3 && edit_y == 8) ? ((X3 + 11 < x && x < X3 + 56) && Y8 + 47 == y) :
                (edit_x == 4 && edit_y == 8) ? ((X4 + 11 < x && x < X4 + 56) && Y8 + 47 == y) :
                (edit_x == 5 && edit_y == 8) ? ((X5 + 11 < x && x < X5 + 56) && Y8 + 47 == y) :
                (edit_x == 6 && edit_y == 8) ? ((X6 + 11 < x && x < X6 + 56) && Y8 + 47 == y) :
                (edit_x == 7 && edit_y == 8) ? ((X7 + 11 < x && x < X7 + 56) && Y8 + 47 == y) :
                (edit_x == 8 && edit_y == 8) ? ((X8 + 11 < x && x < X8 + 56) && Y8 + 47 == y) :
                0;

                
 
 ///////////////////////////number_print/////////////////////////////////////////////////
 assign num[0] = (array[3:0] == 4'b0001) ? (x > X0 + 30 && x < X0 + 42 && y > Y0 + 6 && y < Y0 + 48) :



              (array[3:0] == 4'b0010) ? ((x > X0 + 20 && x < X0 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y0 + 30 && y < Y0 + 42)) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y0 + 42 && y < Y0 + 48):


                
              (array[3:0] == 4'b0011) ? (x > X0 + 20 && x < X0 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y0 + 42 && y < Y0 + 48):

  
              (array[3:0] == 4'b0100) ? (x > X0 + 20 && x < X0 + 27 && y > Y0 + 6 && y < Y0 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y0 + 6 && y < Y0 + 48): 


             (array[3:0] == 4'b0101) ? (x > X0 + 20 && x < X0 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y0 + 42 && y < Y0 + 48) :

             (array[3:0] == 4'b0110) ? (x > X0 + 20 && x < X0 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        
             (array[3:0] == 4'b0111) ?   (x > X0 + 20 && x < X0 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y0 + 12 && y < Y0 + 48) : 


             (array[3:0] == 4'b1000) ? (x > X0 + 20 && x < X0 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X0 + 45 && x < X0 + 52 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                         
             (array[3:0] == 4'b1001) ?  (x > X0 + 20 && x < X0 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                        (x > X0 + 20 && x < X0 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X0 + 45 && x < X0 + 52 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                        (x > X0 + 20 && x < X0 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        0;

assign num[1] = (array[7:4] == 4'b0001) ? (x > X1 + 30 && x < X1 + 42 && y > Y0 + 6 && y < Y0 + 48) :



              (array[7:4] == 4'b0010) ? ((x > X1 + 20 && x < X1 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y0 + 30 && y < Y0 + 42)) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y0 + 42 && y < Y0 + 48):


                
              (array[7:4] == 4'b0011) ? (x > X1 + 20 && x < X1 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y0 + 42 && y < Y0 + 48):

  
              (array[7:4] == 4'b0100) ? (x > X1 + 20 && x < X1 + 27 && y > Y0 + 6 && y < Y0 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y0 + 6 && y < Y0 + 48): 


             (array[7:4] == 4'b0101) ? (x > X1 + 20 && x < X1 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y0 + 42 && y < Y0 + 48) :

             (array[7:4] == 4'b0110) ? (x > X1 + 20 && x < X1 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        
             (array[7:4] == 4'b0111) ?   (x > X1 + 20 && x < X1 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y0 + 12 && y < Y0 + 48) : 


             (array[7:4] == 4'b1000) ? (x > X1 + 20 && x < X1 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X1 + 45 && x < X1 + 52 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                         
             (array[7:4] == 4'b1001) ?  (x > X1 + 20 && x < X1 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                        (x > X1 + 20 && x < X1 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X1 + 45 && x < X1 + 52 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                        (x > X1 + 20 && x < X1 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        0;

assign num[2] = (array[11:8] == 4'b0001) ? (x > X2 + 30 && x < X2 + 42 && y > Y0 + 6 && y < Y0 + 48) :



              (array[11:8] == 4'b0010) ? ((x > X2 + 20 && x < X2 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y0 + 30 && y < Y0 + 42)) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y0 + 42 && y < Y0 + 48):


                
              (array[11:8] == 4'b0011) ? (x > X2 + 20 && x < X2 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y0 + 42 && y < Y0 + 48):

  
              (array[11:8] == 4'b0100) ? (x > X2 + 20 && x < X2 + 27 && y > Y0 + 6 && y < Y0 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y0 + 6 && y < Y0 + 48): 


             (array[11:8] == 4'b0101) ? (x > X2 + 20 && x < X2 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y0 + 42 && y < Y0 + 48) :

             (array[11:8] == 4'b0110) ? (x > X2 + 20 && x < X2 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        
             (array[11:8] == 4'b0111) ?   (x > X2 + 20 && x < X2 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y0 + 12 && y < Y0 + 48) : 


             (array[11:8] == 4'b1000) ? (x > X2 + 20 && x < X2 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X2 + 45 && x < X2 + 52 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                         
             (array[11:8] == 4'b1001) ?  (x > X2 + 20 && x < X2 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                        (x > X2 + 20 && x < X2 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X2 + 45 && x < X2 + 52 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                        (x > X2 + 20 && x < X2 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        0;


assign num[3] = (array[15:12] == 4'b0001) ? (x > X3 + 30 && x < X3 + 42 && y > Y0 + 6 && y < Y0 + 48) :



              (array[15:12] == 4'b0010) ? ((x > X3 + 20 && x < X3 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y0 + 30 && y < Y0 + 42)) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y0 + 42 && y < Y0 + 48):


                
              (array[15:12] == 4'b0011) ? (x > X3 + 20 && x < X3 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y0 + 42 && y < Y0 + 48):

  
              (array[15:12] == 4'b0100) ? (x > X3 + 20 && x < X3 + 27 && y > Y0 + 6 && y < Y0 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y0 + 6 && y < Y0 + 48): 


             (array[15:12] == 4'b0101) ? (x > X3 + 20 && x < X3 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y0 + 42 && y < Y0 + 48) :

             (array[15:12] == 4'b0110) ? (x > X3 + 20 && x < X3 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        
             (array[15:12] == 4'b0111) ?   (x > X3 + 20 && x < X3 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y0 + 12 && y < Y0 + 48) : 


             (array[15:12] == 4'b1000) ? (x > X3 + 20 && x < X3 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X3 + 45 && x < X3 + 52 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                         
             (array[15:12] == 4'b1001) ?  (x > X3 + 20 && x < X3 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                        (x > X3 + 20 && x < X3 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X3 + 45 && x < X3 + 52 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                        (x > X3 + 20 && x < X3 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        0;


assign num[4] = (array[19:16] == 4'b0001) ? (x > X4 + 30 && x < X4 + 42 && y > Y0 + 6 && y < Y0 + 48) :



              (array[19:16] == 4'b0010) ? ((x > X4 + 20 && x < X4 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y0 + 30 && y < Y0 + 42)) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y0 + 42 && y < Y0 + 48):


                
              (array[19:16] == 4'b0011) ? (x > X4 + 20 && x < X4 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y0 + 42 && y < Y0 + 48):

  
              (array[19:16] == 4'b0100) ? (x > X4 + 20 && x < X4 + 27 && y > Y0 + 6 && y < Y0 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y0 + 6 && y < Y0 + 48): 


             (array[19:16] == 4'b0101) ? (x > X4 + 20 && x < X4 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y0 + 42 && y < Y0 + 48) :

             (array[19:16] == 4'b0110) ? (x > X4 + 20 && x < X4 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        
             (array[19:16] == 4'b0111) ?   (x > X4 + 20 && x < X4 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y0 + 12 && y < Y0 + 48) : 


             (array[19:16] == 4'b1000) ? (x > X4 + 20 && x < X4 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X4 + 45 && x < X4 + 52 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                         
             (array[19:16] == 4'b1001) ?  (x > X4 + 20 && x < X4 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                        (x > X4 + 20 && x < X4 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X4 + 45 && x < X4 + 52 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                        (x > X4 + 20 && x < X4 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        0;

assign num[5] = (array[23:20] == 4'b0001) ? (x > X5 + 30 && x < X5 + 42 && y > Y0 + 6 && y < Y0 + 48) :



              (array[23:20] == 4'b0010) ? ((x > X5 + 20 && x < X5 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y0 + 30 && y < Y0 + 42)) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y0 + 42 && y < Y0 + 48):


                
              (array[23:20] == 4'b0011) ? (x > X5 + 20 && x < X5 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y0 + 42 && y < Y0 + 48):

  
              (array[23:20] == 4'b0100) ? (x > X5 + 20 && x < X5 + 27 && y > Y0 + 6 && y < Y0 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y0 + 6 && y < Y0 + 48): 


             (array[23:20] == 4'b0101) ? (x > X5 + 20 && x < X5 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y0 + 42 && y < Y0 + 48) :

             (array[23:20] == 4'b0110) ? (x > X5 + 20 && x < X5 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        
             (array[23:20] == 4'b0111) ?   (x > X5 + 20 && x < X5 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y0 + 12 && y < Y0 + 48) : 


             (array[23:20] == 4'b1000) ? (x > X5 + 20 && x < X5 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X5 + 45 && x < X5 + 52 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                         
             (array[23:20] == 4'b1001) ?  (x > X5 + 20 && x < X5 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                        (x > X5 + 20 && x < X5 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X5 + 45 && x < X5 + 52 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                        (x > X5 + 20 && x < X5 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        0;


assign num[6] = (array[27:24] == 4'b0001) ? (x > X6 + 30 && x < X6 + 42 && y > Y0 + 6 && y < Y0 + 48) :



              (array[27:24] == 4'b0010) ? ((x > X6 + 20 && x < X6 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y0 + 30 && y < Y0 + 42)) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y0 + 42 && y < Y0 + 48):


                
              (array[27:24] == 4'b0011) ? (x > X6 + 20 && x < X6 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y0 + 42 && y < Y0 + 48):

  
              (array[27:24] == 4'b0100) ? (x > X6 + 20 && x < X6 + 27 && y > Y0 + 6 && y < Y0 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y0 + 6 && y < Y0 + 48): 


             (array[27:24] == 4'b0101) ? (x > X6 + 20 && x < X6 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y0 + 42 && y < Y0 + 48) :

             (array[27:24] == 4'b0110) ? (x > X6 + 20 && x < X6 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        
             (array[27:24] == 4'b0111) ?   (x > X6 + 20 && x < X6 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y0 + 12 && y < Y0 + 48) : 


             (array[27:24] == 4'b1000) ? (x > X6 + 20 && x < X6 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X6 + 45 && x < X6 + 52 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                         
             (array[27:24] == 4'b1001) ?  (x > X6 + 20 && x < X6 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                        (x > X6 + 20 && x < X6 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X6 + 45 && x < X6 + 52 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                        (x > X6 + 20 && x < X6 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        0;


assign num[7] = (array[31:28] == 4'b0001) ? (x > X7 + 30 && x < X7 + 42 && y > Y0 + 6 && y < Y0 + 48) :



              (array[31:28] == 4'b0010) ? ((x > X7 + 20 && x < X7 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y0 + 30 && y < Y0 + 42)) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y0 + 42 && y < Y0 + 48):


                
              (array[31:28] == 4'b0011) ? (x > X7 + 20 && x < X7 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y0 + 42 && y < Y0 + 48):

  
              (array[31:28] == 4'b0100) ? (x > X7 + 20 && x < X7 + 27 && y > Y0 + 6 && y < Y0 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y0 + 6 && y < Y0 + 48): 


             (array[31:28] == 4'b0101) ? (x > X7 + 20 && x < X7 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y0 + 42 && y < Y0 + 48) :

             (array[31:28] == 4'b0110) ? (x > X7 + 20 && x < X7 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        
             (array[31:28] == 4'b0111) ?   (x > X7 + 20 && x < X7 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y0 + 12 && y < Y0 + 48) : 


             (array[31:28] == 4'b1000) ? (x > X7 + 20 && x < X7 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X7 + 45 && x < X7 + 52 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                         
             (array[31:28] == 4'b1001) ?  (x > X7 + 20 && x < X7 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                        (x > X7 + 20 && x < X7 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X7 + 45 && x < X7 + 52 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                        (x > X7 + 20 && x < X7 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        0;
assign num[8] = (array[35:32] == 4'b0001) ? (x > X8 + 30 && x < X8 + 42 && y > Y0 + 6 && y < Y0 + 48) :



              (array[35:32] == 4'b0010) ? ((x > X8 + 20 && x < X8 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y0 + 30 && y < Y0 + 42)) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y0 + 42 && y < Y0 + 48):


                
              (array[35:32] == 4'b0011) ? (x > X8 + 20 && x < X8 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y0 + 12 && y < Y0 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y0 + 42 && y < Y0 + 48):

  
              (array[35:32] == 4'b0100) ? (x > X8 + 20 && x < X8 + 27 && y > Y0 + 6 && y < Y0 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y0 + 6 && y < Y0 + 48): 


             (array[35:32] == 4'b0101) ? (x > X8 + 20 && x < X8 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y0 + 42 && y < Y0 + 48) :

             (array[35:32] == 4'b0110) ? (x > X8 + 20 && x < X8 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y0 + 24 && y < Y0 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y0 + 30 && y < Y0 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        
             (array[35:32] == 4'b0111) ?   (x > X8 + 20 && x < X8 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y0 + 12 && y < Y0 + 48) : 


             (array[35:32] == 4'b1000) ? (x > X8 + 20 && x < X8 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X8 + 45 && x < X8 + 52 && y > Y0 + 12 && y < Y0 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                         
             (array[35:32] == 4'b1001) ?  (x > X8 + 20 && x < X8 + 52 && y > Y0 + 6 && y < Y0 + 12) || 
                                        (x > X8 + 20 && x < X8 + 27 && y > Y0 + 12 && y < Y0 + 24) || 
                                        (x > X8 + 45 && x < X8 + 52 && y > Y0 + 12 && y < Y0 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y0 + 24 && y < Y0 + 30) ||
                                        (x > X8 + 20 && x < X8 + 52 && y > Y0 + 42 && y < Y0 + 48) : 
                                        0;
////////////////////////////////////////line2///////////////////////////////////////////////////////////////////////                
                assign num[9] = (array[39:36] == 4'b0001) ? (x > X0 + 30 && x < X0 + 42 && y > Y1 + 6 && y < Y1 + 48) :



              (array[39:36] == 4'b0010) ? ((x > X0 + 20 && x < X0 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y1 + 30 && y < Y1 + 42)) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y1 + 42 && y < Y1 + 48):


                
              (array[39:36] == 4'b0011) ? (x > X0 + 20 && x < X0 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y1 + 42 && y < Y1 + 48):

  
              (array[39:36] == 4'b0100) ? (x > X0 + 20 && x < X0 + 27 && y > Y1 + 6 && y < Y1 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y1 + 6 && y < Y1 + 48): 


             (array[39:36] == 4'b0101) ? (x > X0 + 20 && x < X0 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y1 + 42 && y < Y1 + 48) :

             (array[39:36] == 4'b0110) ? (x > X0 + 20 && x < X0 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        
             (array[39:36] == 4'b0111) ?   (x > X0 + 20 && x < X0 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y1 + 12 && y < Y1 + 48) : 


             (array[39:36] == 4'b1000) ? (x > X0 + 20 && x < X0 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X0 + 45 && x < X0 + 52 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                         
             (array[39:36] == 4'b1001) ?  (x > X0 + 20 && x < X0 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                        (x > X0 + 20 && x < X0 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X0 + 45 && x < X0 + 52 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                        (x > X0 + 20 && x < X0 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        0;

assign num[10] = (array[43:40] == 4'b0001) ? (x > X1 + 30 && x < X1 + 42 && y > Y1 + 6 && y < Y1 + 48) :



              (array[43:40] == 4'b0010) ? ((x > X1 + 20 && x < X1 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y1 + 30 && y < Y1 + 42)) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y1 + 42 && y < Y1 + 48):


                
              (array[43:40] == 4'b0011) ? (x > X1 + 20 && x < X1 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y1 + 42 && y < Y1 + 48):

  
              (array[43:40] == 4'b0100) ? (x > X1 + 20 && x < X1 + 27 && y > Y1 + 6 && y < Y1 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y1 + 6 && y < Y1 + 48): 


             (array[43:40] == 4'b0101) ? (x > X1 + 20 && x < X1 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y1 + 42 && y < Y1 + 48) :

             (array[43:40] == 4'b0110) ? (x > X1 + 20 && x < X1 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        
             (array[43:40] == 4'b0111) ?   (x > X1 + 20 && x < X1 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y1 + 12 && y < Y1 + 48) : 


             (array[43:40] == 4'b1000) ? (x > X1 + 20 && x < X1 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X1 + 45 && x < X1 + 52 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                         
             (array[43:40] == 4'b1001) ?  (x > X1 + 20 && x < X1 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                        (x > X1 + 20 && x < X1 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X1 + 45 && x < X1 + 52 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                        (x > X1 + 20 && x < X1 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        0;

assign num[11] = (array[47:44] == 4'b0001) ? (x > X2 + 30 && x < X2 + 42 && y > Y1 + 6 && y < Y1 + 48) :



              (array[47:44] == 4'b0010) ? ((x > X2 + 20 && x < X2 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y1 + 30 && y < Y1 + 42)) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y1 + 42 && y < Y1 + 48):


                
              (array[47:44] == 4'b0011) ? (x > X2 + 20 && x < X2 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y1 + 42 && y < Y1 + 48):

  
              (array[47:44] == 4'b0100) ? (x > X2 + 20 && x < X2 + 27 && y > Y1 + 6 && y < Y1 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y1 + 6 && y < Y1 + 48): 


             (array[47:44] == 4'b0101) ? (x > X2 + 20 && x < X2 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y1 + 42 && y < Y1 + 48) :

             (array[47:44] == 4'b0110) ? (x > X2 + 20 && x < X2 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        
             (array[47:44] == 4'b0111) ?   (x > X2 + 20 && x < X2 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y1 + 12 && y < Y1 + 48) : 


             (array[47:44] == 4'b1000) ? (x > X2 + 20 && x < X2 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X2 + 45 && x < X2 + 52 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                         
             (array[47:44] == 4'b1001) ?  (x > X2 + 20 && x < X2 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                        (x > X2 + 20 && x < X2 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X2 + 45 && x < X2 + 52 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                        (x > X2 + 20 && x < X2 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        0;
assign num[12] = (array[51:48] == 4'b0001) ? (x > X3 + 30 && x < X3 + 42 && y > Y1 + 6 && y < Y1 + 48) :



              (array[51:48] == 4'b0010) ? ((x > X3 + 20 && x < X3 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y1 + 30 && y < Y1 + 42)) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y1 + 42 && y < Y1 + 48):


                
              (array[51:48] == 4'b0011) ? (x > X3 + 20 && x < X3 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y1 + 42 && y < Y1 + 48):

  
              (array[51:48] == 4'b0100) ? (x > X3 + 20 && x < X3 + 27 && y > Y1 + 6 && y < Y1 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y1 + 6 && y < Y1 + 48): 


             (array[51:48] == 4'b0101) ? (x > X3 + 20 && x < X3 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y1 + 42 && y < Y1 + 48) :

             (array[51:48] == 4'b0110) ? (x > X3 + 20 && x < X3 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        
             (array[51:48] == 4'b0111) ?   (x > X3 + 20 && x < X3 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y1 + 12 && y < Y1 + 48) : 


             (array[51:48] == 4'b1000) ? (x > X3 + 20 && x < X3 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X3 + 45 && x < X3 + 52 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                         
             (array[51:48] == 4'b1001) ?  (x > X3 + 20 && x < X3 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                        (x > X3 + 20 && x < X3 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X3 + 45 && x < X3 + 52 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                        (x > X3 + 20 && x < X3 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        0;

assign num[13] = (array[55:52] == 4'b0001) ? (x > X4 + 30 && x < X4 + 42 && y > Y1 + 6 && y < Y1 + 48) :



              (array[55:52] == 4'b0010) ? ((x > X4 + 20 && x < X4 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y1 + 30 && y < Y1 + 42)) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y1 + 42 && y < Y1 + 48):


                
              (array[55:52] == 4'b0011) ? (x > X4 + 20 && x < X4 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y1 + 42 && y < Y1 + 48):

  
              (array[55:52] == 4'b0100) ? (x > X4 + 20 && x < X4 + 27 && y > Y1 + 6 && y < Y1 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y1 + 6 && y < Y1 + 48): 


             (array[55:52] == 4'b0101) ? (x > X4 + 20 && x < X4 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y1 + 42 && y < Y1 + 48) :

             (array[55:52] == 4'b0110) ? (x > X4 + 20 && x < X4 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        
             (array[55:52] == 4'b0111) ?   (x > X4 + 20 && x < X4 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y1 + 12 && y < Y1 + 48) : 


             (array[55:52] == 4'b1000) ? (x > X4 + 20 && x < X4 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X4 + 45 && x < X4 + 52 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                         
             (array[55:52] == 4'b1001) ?  (x > X4 + 20 && x < X4 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                        (x > X4 + 20 && x < X4 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X4 + 45 && x < X4 + 52 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                        (x > X4 + 20 && x < X4 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        0;

assign num[14] = (array[59:56] == 4'b0001) ? (x > X5 + 30 && x < X5 + 42 && y > Y1 + 6 && y < Y1 + 48) :



              (array[59:56] == 4'b0010) ? ((x > X5 + 20 && x < X5 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y1 + 30 && y < Y1 + 42)) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y1 + 42 && y < Y1 + 48):


                
              (array[59:56] == 4'b0011) ? (x > X5 + 20 && x < X5 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y1 + 42 && y < Y1 + 48):

  
              (array[59:56] == 4'b0100) ? (x > X5 + 20 && x < X5 + 27 && y > Y1 + 6 && y < Y1 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y1 + 6 && y < Y1 + 48): 


             (array[59:56] == 4'b0101) ? (x > X5 + 20 && x < X5 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y1 + 42 && y < Y1 + 48) :

             (array[59:56] == 4'b0110) ? (x > X5 + 20 && x < X5 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        
             (array[59:56] == 4'b0111) ?   (x > X5 + 20 && x < X5 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y1 + 12 && y < Y1 + 48) : 


             (array[59:56] == 4'b1000) ? (x > X5 + 20 && x < X5 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X5 + 45 && x < X5 + 52 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                         
             (array[59:56] == 4'b1001) ?  (x > X5 + 20 && x < X5 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                        (x > X5 + 20 && x < X5 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X5 + 45 && x < X5 + 52 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                        (x > X5 + 20 && x < X5 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        0;

assign num[15] = (array[63:60] == 4'b0001) ? (x > X6 + 30 && x < X6 + 42 && y > Y1 + 6 && y < Y1 + 48) :



              (array[63:60] == 4'b0010) ? ((x > X6 + 20 && x < X6 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y1 + 30 && y < Y1 + 42)) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y1 + 42 && y < Y1 + 48):


                
              (array[63:60] == 4'b0011) ? (x > X6 + 20 && x < X6 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y1 + 42 && y < Y1 + 48):

  
              (array[63:60] == 4'b0100) ? (x > X6 + 20 && x < X6 + 27 && y > Y1 + 6 && y < Y1 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y1 + 6 && y < Y1 + 48): 


             (array[63:60] == 4'b0101) ? (x > X6 + 20 && x < X6 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y1 + 42 && y < Y1 + 48) :

             (array[63:60] == 4'b0110) ? (x > X6 + 20 && x < X6 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        
             (array[63:60] == 4'b0111) ?   (x > X6 + 20 && x < X6 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y1 + 12 && y < Y1 + 48) : 


             (array[63:60] == 4'b1000) ? (x > X6 + 20 && x < X6 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X6 + 45 && x < X6 + 52 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                         
             (array[63:60] == 4'b1001) ?  (x > X6 + 20 && x < X6 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                        (x > X6 + 20 && x < X6 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X6 + 45 && x < X6 + 52 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                        (x > X6 + 20 && x < X6 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        0;
assign num[16] = (array[67:64] == 4'b0001) ? (x > X7 + 30 && x < X7 + 42 && y > Y1 + 6 && y < Y1 + 48) :



              (array[67:64] == 4'b0010) ? ((x > X7 + 20 && x < X7 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y1 + 30 && y < Y1 + 42)) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y1 + 42 && y < Y1 + 48):


                
              (array[67:64] == 4'b0011) ? (x > X7 + 20 && x < X7 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y1 + 42 && y < Y1 + 48):

  
              (array[67:64] == 4'b0100) ? (x > X7 + 20 && x < X7 + 27 && y > Y1 + 6 && y < Y1 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y1 + 6 && y < Y1 + 48): 


             (array[67:64] == 4'b0101) ? (x > X7 + 20 && x < X7 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y1 + 42 && y < Y1 + 48) :

             (array[67:64] == 4'b0110) ? (x > X7 + 20 && x < X7 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        
             (array[67:64] == 4'b0111) ?   (x > X7 + 20 && x < X7 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y1 + 12 && y < Y1 + 48) : 


             (array[67:64] == 4'b1000) ? (x > X7 + 20 && x < X7 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X7 + 45 && x < X7 + 52 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                         
             (array[67:64] == 4'b1001) ?  (x > X7 + 20 && x < X7 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                        (x > X7 + 20 && x < X7 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X7 + 45 && x < X7 + 52 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                        (x > X7 + 20 && x < X7 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        0;

assign num[17] = (array[71:68] == 4'b0001) ? (x > X8 + 30 && x < X8 + 42 && y > Y1 + 6 && y < Y1 + 48) :



              (array[71:68] == 4'b0010) ? ((x > X8 + 20 && x < X8 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y1 + 30 && y < Y1 + 42)) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y1 + 42 && y < Y1 + 48):


                
              (array[71:68] == 4'b0011) ? (x > X8 + 20 && x < X8 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y1 + 12 && y < Y1 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y1 + 42 && y < Y1 + 48):

  
              (array[71:68] == 4'b0100) ? (x > X8 + 20 && x < X8 + 27 && y > Y1 + 6 && y < Y1 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y1 + 6 && y < Y1 + 48): 


             (array[71:68] == 4'b0101) ? (x > X8 + 20 && x < X8 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y1 + 42 && y < Y1 + 48) :

             (array[71:68] == 4'b0110) ? (x > X8 + 20 && x < X8 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y1 + 24 && y < Y1 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y1 + 30 && y < Y1 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        
             (array[71:68] == 4'b0111) ?   (x > X8 + 20 && x < X8 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y1 + 12 && y < Y1 + 48) : 


             (array[71:68] == 4'b1000) ? (x > X8 + 20 && x < X8 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X8 + 45 && x < X8 + 52 && y > Y1 + 12 && y < Y1 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                         
             (array[71:68] == 4'b1001) ?  (x > X8 + 20 && x < X8 + 52 && y > Y1 + 6 && y < Y1 + 12) || 
                                        (x > X8 + 20 && x < X8 + 27 && y > Y1 + 12 && y < Y1 + 24) || 
                                        (x > X8 + 45 && x < X8 + 52 && y > Y1 + 12 && y < Y1 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y1 + 24 && y < Y1 + 30) ||
                                        (x > X8 + 20 && x < X8 + 52 && y > Y1 + 42 && y < Y1 + 48) : 
                                        0;
                                        
                                        
  //////////////////////////////////////////////////line3////////////////////////////////////////////////////
          assign num[18] = (array[75:72] == 4'b0001) ? (x > X0 + 30 && x < X0 + 42 && y > Y2 + 6 && y < Y2 + 48) :



              (array[75:72] == 4'b0010) ? ((x > X0 + 20 && x < X0 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y2 + 30 && y < Y2 + 42)) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y2 + 42 && y < Y2 + 48):

                
              (array[75:72] == 4'b0011) ? (x > X0 + 20 && x < X0 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y2 + 42 && y < Y2 + 48):

  
              (array[75:72] == 4'b0100) ? (x > X0 + 20 && x < X0 + 27 && y > Y2 + 6 && y < Y2 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y2 + 6 && y < Y2 + 48): 


             (array[75:72] == 4'b0101) ? (x > X0 + 20 && x < X0 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y2 + 42 && y < Y2 + 48) :

             (array[75:72] == 4'b0110) ? (x > X0 + 20 && x < X0 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        
             (array[75:72] == 4'b0111) ?   (x > X0 + 20 && x < X0 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y2 + 12 && y < Y2 + 48) : 


             (array[75:72] == 4'b1000) ? (x > X0 + 20 && x < X0 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X0 + 45 && x < X0 + 52 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                         
             (array[75:72] == 4'b1001) ?  (x > X0 + 20 && x < X0 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                        (x > X0 + 20 && x < X0 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X0 + 45 && x < X0 + 52 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                        (x > X0 + 20 && x < X0 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        0;      
                





        assign num[19] = (array[79:76] == 4'b0001) ? (x > X1 + 30 && x < X1 + 42 && y > Y2 + 6 && y < Y2 + 48) :



              (array[79:76] == 4'b0010) ? ((x > X1 + 20 && x < X1 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y2 + 30 && y < Y2 + 42)) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y2 + 42 && y < Y2 + 48):

                
              (array[79:76] == 4'b0011) ? (x > X1 + 20 && x < X1 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y2 + 42 && y < Y2 + 48):

  
              (array[79:76] == 4'b0100) ? (x > X1 + 20 && x < X1 + 27 && y > Y2 + 6 && y < Y2 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y2 + 6 && y < Y2 + 48): 


             (array[79:76] == 4'b0101) ? (x > X1 + 20 && x < X1 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y2 + 42 && y < Y2 + 48) :

             (array[79:76] == 4'b0110) ? (x > X1 + 20 && x < X1 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        
             (array[79:76] == 4'b0111) ?   (x > X1 + 20 && x < X1 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y2 + 12 && y < Y2 + 48) : 


             (array[79:76] == 4'b1000) ? (x > X1 + 20 && x < X1 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X1 + 45 && x < X1 + 52 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                         
             (array[79:76] == 4'b1001) ?  (x > X1 + 20 && x < X1 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                        (x > X1 + 20 && x < X1 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X1 + 45 && x < X1 + 52 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                        (x > X1 + 20 && x < X1 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        0;      
                
  


        assign num[20] = (array[83:80] == 4'b0001) ? (x > X2 + 30 && x < X2 + 42 && y > Y2 + 6 && y < Y2 + 48) :



              (array[83:80] == 4'b0010) ? ((x > X2 + 20 && x < X2 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y2 + 30 && y < Y2 + 42)) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y2 + 42 && y < Y2 + 48):

                
              (array[83:80] == 4'b0011) ? (x > X2 + 20 && x < X2 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y2 + 42 && y < Y2 + 48):

  
              (array[83:80] == 4'b0100) ? (x > X2 + 20 && x < X2 + 27 && y > Y2 + 6 && y < Y2 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y2 + 6 && y < Y2 + 48): 


             (array[83:80] == 4'b0101) ? (x > X2 + 20 && x < X2 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y2 + 42 && y < Y2 + 48) :

             (array[83:80] == 4'b0110) ? (x > X2 + 20 && x < X2 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        
             (array[83:80] == 4'b0111) ?   (x > X2 + 20 && x < X2 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y2 + 12 && y < Y2 + 48) : 


             (array[83:80] == 4'b1000) ? (x > X2 + 20 && x < X2 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X2 + 45 && x < X2 + 52 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                         
             (array[83:80] == 4'b1001) ?  (x > X2 + 20 && x < X2 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                        (x > X2 + 20 && x < X2 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X2 + 45 && x < X2 + 52 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                        (x > X2 + 20 && x < X2 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        0;      



        assign num[21] = (array[87:84] == 4'b0001) ? (x > X3 + 30 && x < X3 + 42 && y > Y2 + 6 && y < Y2 + 48) :



              (array[87:84] == 4'b0010) ? ((x > X3 + 20 && x < X3 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y2 + 30 && y < Y2 + 42)) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y2 + 42 && y < Y2 + 48):

                
              (array[87:84] == 4'b0011) ? (x > X3 + 20 && x < X3 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y2 + 42 && y < Y2 + 48):

  
              (array[87:84] == 4'b0100) ? (x > X3 + 20 && x < X3 + 27 && y > Y2 + 6 && y < Y2 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y2 + 6 && y < Y2 + 48): 


             (array[87:84] == 4'b0101) ? (x > X3 + 20 && x < X3 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y2 + 42 && y < Y2 + 48) :

             (array[87:84] == 4'b0110) ? (x > X3 + 20 && x < X3 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        
             (array[87:84] == 4'b0111) ?   (x > X3 + 20 && x < X3 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y2 + 12 && y < Y2 + 48) : 


             (array[87:84] == 4'b1000) ? (x > X3 + 20 && x < X3 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X3 + 45 && x < X3 + 52 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                         
             (array[87:84] == 4'b1001) ?  (x > X3 + 20 && x < X3 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                        (x > X3 + 20 && x < X3 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X3 + 45 && x < X3 + 52 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                        (x > X3 + 20 && x < X3 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        0;      
                
  



        assign num[22] = (array[91:88] == 4'b0001) ? (x > X4 + 30 && x < X4 + 42 && y > Y2 + 6 && y < Y2 + 48) :



              (array[91:88] == 4'b0010) ? ((x > X4 + 20 && x < X4 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y2 + 30 && y < Y2 + 42)) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y2 + 42 && y < Y2 + 48):

                
              (array[91:88] == 4'b0011) ? (x > X4 + 20 && x < X4 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y2 + 42 && y < Y2 + 48):

  
              (array[91:88] == 4'b0100) ? (x > X4 + 20 && x < X4 + 27 && y > Y2 + 6 && y < Y2 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y2 + 6 && y < Y2 + 48): 


             (array[91:88] == 4'b0101) ? (x > X4 + 20 && x < X4 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y2 + 42 && y < Y2 + 48) :

             (array[91:88] == 4'b0110) ? (x > X4 + 20 && x < X4 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        
             (array[91:88] == 4'b0111) ?   (x > X4 + 20 && x < X4 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y2 + 12 && y < Y2 + 48) : 


             (array[91:88] == 4'b1000) ? (x > X4 + 20 && x < X4 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X4 + 45 && x < X4 + 52 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                         
             (array[91:88] == 4'b1001) ?  (x > X4 + 20 && x < X4 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                        (x > X4 + 20 && x < X4 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X4 + 45 && x < X4 + 52 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                        (x > X4 + 20 && x < X4 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        0;      
                
  
                
  
          assign num[23] = (array[95:92] == 4'b0001) ? (x > X5 + 30 && x < X5 + 42 && y > Y2 + 6 && y < Y2 + 48) :



              (array[95:92] == 4'b0010) ? ((x > X5 + 20 && x < X5 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y2 + 30 && y < Y2 + 42)) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y2 + 42 && y < Y2 + 48):

                
              (array[95:92] == 4'b0011) ? (x > X5 + 20 && x < X5 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y2 + 42 && y < Y2 + 48):

  
              (array[95:92] == 4'b0100) ? (x > X5 + 20 && x < X5 + 27 && y > Y2 + 6 && y < Y2 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y2 + 6 && y < Y2 + 48): 


             (array[95:92] == 4'b0101) ? (x > X5 + 20 && x < X5 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y2 + 42 && y < Y2 + 48) :

             (array[95:92] == 4'b0110) ? (x > X5 + 20 && x < X5 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        
             (array[95:92] == 4'b0111) ?   (x > X5 + 20 && x < X5 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y2 + 12 && y < Y2 + 48) : 


             (array[95:92] == 4'b1000) ? (x > X5 + 20 && x < X5 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X5 + 45 && x < X5 + 52 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                         
             (array[95:92] == 4'b1001) ?  (x > X5 + 20 && x < X5 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                        (x > X5 + 20 && x < X5 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X5 + 45 && x < X5 + 52 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                        (x > X5 + 20 && x < X5 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        0;      
                
  

        assign num[24] = (array[99:96] == 4'b0001) ? (x > X6 + 30 && x < X6 + 42 && y > Y2 + 6 && y < Y2 + 48) :



              (array[99:96] == 4'b0010) ? ((x > X6 + 20 && x < X6 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y2 + 30 && y < Y2 + 42)) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y2 + 42 && y < Y2 + 48):

                
              (array[99:96] == 4'b0011) ? (x > X6 + 20 && x < X6 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y2 + 42 && y < Y2 + 48):

  
              (array[99:96] == 4'b0100) ? (x > X6 + 20 && x < X6 + 27 && y > Y2 + 6 && y < Y2 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y2 + 6 && y < Y2 + 48): 


             (array[99:96] == 4'b0101) ? (x > X6 + 20 && x < X6 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y2 + 42 && y < Y2 + 48) :

             (array[99:96] == 4'b0110) ? (x > X6 + 20 && x < X6 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        
             (array[99:96] == 4'b0111) ?   (x > X6 + 20 && x < X6 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y2 + 12 && y < Y2 + 48) : 


             (array[99:96] == 4'b1000) ? (x > X6 + 20 && x < X6 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X6 + 45 && x < X6 + 52 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                         
             (array[99:96] == 4'b1001) ?  (x > X6 + 20 && x < X6 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                        (x > X6 + 20 && x < X6 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X6 + 45 && x < X6 + 52 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                        (x > X6 + 20 && x < X6 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        0;      
                
  
        assign num[25] = (array[103:100] == 4'b0001) ? (x > X7 + 30 && x < X7 + 42 && y > Y2 + 6 && y < Y2 + 48) :



              (array[103:100] == 4'b0010) ? ((x > X7 + 20 && x < X7 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y2 + 30 && y < Y2 + 42)) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y2 + 42 && y < Y2 + 48):

                
              (array[103:100] == 4'b0011) ? (x > X7 + 20 && x < X7 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y2 + 42 && y < Y2 + 48):

  
              (array[103:100] == 4'b0100) ? (x > X7 + 20 && x < X7 + 27 && y > Y2 + 6 && y < Y2 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y2 + 6 && y < Y2 + 48): 


             (array[103:100] == 4'b0101) ? (x > X7 + 20 && x < X7 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y2 + 42 && y < Y2 + 48) :

             (array[103:100] == 4'b0110) ? (x > X7 + 20 && x < X7 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        
             (array[103:100] == 4'b0111) ?   (x > X7 + 20 && x < X7 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y2 + 12 && y < Y2 + 48) : 


             (array[103:100] == 4'b1000) ? (x > X7 + 20 && x < X7 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X7 + 45 && x < X7 + 52 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                         
             (array[103:100] == 4'b1001) ?  (x > X7 + 20 && x < X7 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                        (x > X7 + 20 && x < X7 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X7 + 45 && x < X7 + 52 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                        (x > X7 + 20 && x < X7 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        0;    



        assign num[26] = (array[107:104] == 4'b0001) ? (x > X8 + 30 && x < X8 + 42 && y > Y2 + 6 && y < Y2 + 48) :



              (array[107:104] == 4'b0010) ? ((x > X8 + 20 && x < X8 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y2 + 30 && y < Y2 + 42)) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y2 + 42 && y < Y2 + 48):

                
              (array[107:104] == 4'b0011) ? (x > X8 + 20 && x < X8 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y2 + 12 && y < Y2 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y2 + 42 && y < Y2 + 48):

  
              (array[107:104] == 4'b0100) ? (x > X8 + 20 && x < X8 + 27 && y > Y2 + 6 && y < Y2 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y2 + 6 && y < Y2 + 48): 


             (array[107:104] == 4'b0101) ? (x > X8 + 20 && x < X8 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y2 + 42 && y < Y2 + 48) :

             (array[107:104] == 4'b0110) ? (x > X8 + 20 && x < X8 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y2 + 24 && y < Y2 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y2 + 30 && y < Y2 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        
             (array[107:104] == 4'b0111) ?   (x > X8 + 20 && x < X8 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y2 + 12 && y < Y2 + 48) : 


             (array[107:104] == 4'b1000) ? (x > X8 + 20 && x < X8 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X8 + 45 && x < X8 + 52 && y > Y2 + 12 && y < Y2 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                         
             (array[107:104] == 4'b1001) ?  (x > X8 + 20 && x < X8 + 52 && y > Y2 + 6 && y < Y2 + 12) || 
                                        (x > X8 + 20 && x < X8 + 27 && y > Y2 + 12 && y < Y2 + 24) || 
                                        (x > X8 + 45 && x < X8 + 52 && y > Y2 + 12 && y < Y2 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y2 + 24 && y < Y2 + 30) ||
                                        (x > X8 + 20 && x < X8 + 52 && y > Y2 + 42 && y < Y2 + 48) : 
                                        0;      
                
    
     ////////////////////////////line4/////////////////////////////////////////////////////////////////
  assign num[27] = (array[111:108] == 4'b0001) ? (x > X0 + 30 && x < X0 + 42 && y > Y3 + 6 && y < Y3 + 48) :



              (array[111:108] == 4'b0010) ? ((x > X0 + 20 && x < X0 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y3 + 30 && y < Y3 + 42)) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y3 + 42 && y < Y3 + 48):


                
              (array[111:108] == 4'b0011) ? (x > X0 + 20 && x < X0 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y3 + 42 && y < Y3 + 48):

  
              (array[111:108] == 4'b0100) ? (x > X0 + 20 && x < X0 + 27 && y > Y3 + 6 && y < Y3 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y3 + 6 && y < Y3 + 48): 


             (array[111:108] == 4'b0101) ? (x > X0 + 20 && x < X0 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y3 + 42 && y < Y3 + 48) :

             (array[111:108] == 4'b0110) ? (x > X0 + 20 && x < X0 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        
             (array[111:108] == 4'b0111) ?   (x > X0 + 20 && x < X0 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y3 + 12 && y < Y3 + 48) : 


             (array[111:108] == 4'b1000) ? (x > X0 + 20 && x < X0 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X0 + 45 && x < X0 + 52 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                         
             (array[111:108] == 4'b1001) ?  (x > X0 + 20 && x < X0 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                        (x > X0 + 20 && x < X0 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X0 + 45 && x < X0 + 52 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                        (x > X0 + 20 && x < X0 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        0;

assign num[28] = (array[115:112] == 4'b0001) ? (x > X1 + 30 && x < X1 + 42 && y > Y3 + 6 && y < Y3 + 48) :



              (array[115:112] == 4'b0010) ? ((x > X1 + 20 && x < X1 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y3 + 30 && y < Y3 + 42)) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y3 + 42 && y < Y3 + 48):


                
              (array[115:112] == 4'b0011) ? (x > X1 + 20 && x < X1 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y3 + 42 && y < Y3 + 48):

  
              (array[115:112] == 4'b0100) ? (x > X1 + 20 && x < X1 + 27 && y > Y3 + 6 && y < Y3 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y3 + 6 && y < Y3 + 48): 


             (array[115:112] == 4'b0101) ? (x > X1 + 20 && x < X1 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y3 + 42 && y < Y3 + 48) :

             (array[115:112] == 4'b0110) ? (x > X1 + 20 && x < X1 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        
             (array[115:112] == 4'b0111) ?   (x > X1 + 20 && x < X1 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y3 + 12 && y < Y3 + 48) : 


             (array[115:112] == 4'b1000) ? (x > X1 + 20 && x < X1 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X1 + 45 && x < X1 + 52 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                         
             (array[115:112] == 4'b1001) ?  (x > X1 + 20 && x < X1 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                        (x > X1 + 20 && x < X1 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X1 + 45 && x < X1 + 52 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                        (x > X1 + 20 && x < X1 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        0;

assign num[29] = (array[119:116] == 4'b0001) ? (x > X2 + 30 && x < X2 + 42 && y > Y3 + 6 && y < Y3 + 48) :



              (array[119:116] == 4'b0010) ? ((x > X2 + 20 && x < X2 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y3 + 30 && y < Y3 + 42)) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y3 + 42 && y < Y3 + 48):


                
              (array[119:116] == 4'b0011) ? (x > X2 + 20 && x < X2 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y3 + 42 && y < Y3 + 48):

  
              (array[119:116] == 4'b0100) ? (x > X2 + 20 && x < X2 + 27 && y > Y3 + 6 && y < Y3 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y3 + 6 && y < Y3 + 48): 


             (array[119:116] == 4'b0101) ? (x > X2 + 20 && x < X2 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y3 + 42 && y < Y3 + 48) :

             (array[119:116] == 4'b0110) ? (x > X2 + 20 && x < X2 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        
             (array[119:116] == 4'b0111) ?   (x > X2 + 20 && x < X2 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y3 + 12 && y < Y3 + 48) : 


             (array[119:116] == 4'b1000) ? (x > X2 + 20 && x < X2 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X2 + 45 && x < X2 + 52 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                         
             (array[119:116] == 4'b1001) ?  (x > X2 + 20 && x < X2 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                        (x > X2 + 20 && x < X2 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X2 + 45 && x < X2 + 52 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                        (x > X2 + 20 && x < X2 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        0;

assign num[30] = (array[123:120] == 4'b0001) ? (x > X3 + 30 && x < X3 + 42 && y > Y3 + 6 && y < Y3 + 48) :



              (array[123:120] == 4'b0010) ? ((x > X3 + 20 && x < X3 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y3 + 30 && y < Y3 + 42)) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y3 + 42 && y < Y3 + 48):


                
              (array[123:120] == 4'b0011) ? (x > X3 + 20 && x < X3 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y3 + 42 && y < Y3 + 48):

  
              (array[123:120] == 4'b0100) ? (x > X3 + 20 && x < X3 + 27 && y > Y3 + 6 && y < Y3 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y3 + 6 && y < Y3 + 48): 


             (array[123:120] == 4'b0101) ? (x > X3 + 20 && x < X3 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y3 + 42 && y < Y3 + 48) :

             (array[123:120] == 4'b0110) ? (x > X3 + 20 && x < X3 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        
             (array[123:120] == 4'b0111) ?   (x > X3 + 20 && x < X3 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y3 + 12 && y < Y3 + 48) : 


             (array[123:120] == 4'b1000) ? (x > X3 + 20 && x < X3 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X3 + 45 && x < X3 + 52 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                         
             (array[123:120] == 4'b1001) ?  (x > X3 + 20 && x < X3 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                        (x > X3 + 20 && x < X3 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X3 + 45 && x < X3 + 52 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                        (x > X3 + 20 && x < X3 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        0;

assign num[31] = (array[127:124] == 4'b0001) ? (x > X4 + 30 && x < X4 + 42 && y > Y3 + 6 && y < Y3 + 48) :



              (array[127:124] == 4'b0010) ? ((x > X4 + 20 && x < X4 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y3 + 30 && y < Y3 + 42)) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y3 + 42 && y < Y3 + 48):


                
              (array[127:124] == 4'b0011) ? (x > X4 + 20 && x < X4 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y3 + 42 && y < Y3 + 48):

  
              (array[127:124] == 4'b0100) ? (x > X4 + 20 && x < X4 + 27 && y > Y3 + 6 && y < Y3 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y3 + 6 && y < Y3 + 48): 


             (array[127:124] == 4'b0101) ? (x > X4 + 20 && x < X4 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y3 + 42 && y < Y3 + 48) :

             (array[127:124] == 4'b0110) ? (x > X4 + 20 && x < X4 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        
             (array[127:124] == 4'b0111) ?   (x > X4 + 20 && x < X4 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y3 + 12 && y < Y3 + 48) : 


             (array[127:124] == 4'b1000) ? (x > X4 + 20 && x < X4 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X4 + 45 && x < X4 + 52 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                         
             (array[127:124] == 4'b1001) ?  (x > X4 + 20 && x < X4 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                        (x > X4 + 20 && x < X4 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X4 + 45 && x < X4 + 52 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                        (x > X4 + 20 && x < X4 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        0;

assign num[32] = (array[131:128] == 4'b0001) ? (x > X5 + 30 && x < X5 + 42 && y > Y3 + 6 && y < Y3 + 48) :



              (array[131:128] == 4'b0010) ? ((x > X5 + 20 && x < X5 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y3 + 30 && y < Y3 + 42)) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y3 + 42 && y < Y3 + 48):


                
              (array[131:128] == 4'b0011) ? (x > X5 + 20 && x < X5 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y3 + 42 && y < Y3 + 48):

  
              (array[131:128] == 4'b0100) ? (x > X5 + 20 && x < X5 + 27 && y > Y3 + 6 && y < Y3 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y3 + 6 && y < Y3 + 48): 


             (array[131:128] == 4'b0101) ? (x > X5 + 20 && x < X5 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y3 + 42 && y < Y3 + 48) :

             (array[131:128] == 4'b0110) ? (x > X5 + 20 && x < X5 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        
             (array[131:128] == 4'b0111) ?   (x > X5 + 20 && x < X5 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y3 + 12 && y < Y3 + 48) : 


             (array[131:128] == 4'b1000) ? (x > X5 + 20 && x < X5 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X5 + 45 && x < X5 + 52 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                         
             (array[131:128] == 4'b1001) ?  (x > X5 + 20 && x < X5 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                        (x > X5 + 20 && x < X5 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X5 + 45 && x < X5 + 52 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                        (x > X5 + 20 && x < X5 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        0;

assign num[33] = (array[135:132] == 4'b0001) ? (x > X6 + 30 && x < X6 + 42 && y > Y3 + 6 && y < Y3 + 48) :



              (array[135:132] == 4'b0010) ? ((x > X6 + 20 && x < X6 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y3 + 30 && y < Y3 + 42)) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y3 + 42 && y < Y3 + 48):


                
              (array[135:132] == 4'b0011) ? (x > X6 + 20 && x < X6 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y3 + 42 && y < Y3 + 48):

  
              (array[135:132] == 4'b0100) ? (x > X6 + 20 && x < X6 + 27 && y > Y3 + 6 && y < Y3 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y3 + 6 && y < Y3 + 48): 


             (array[135:132] == 4'b0101) ? (x > X6 + 20 && x < X6 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y3 + 42 && y < Y3 + 48) :

             (array[135:132] == 4'b0110) ? (x > X6 + 20 && x < X6 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        
             (array[135:132] == 4'b0111) ?   (x > X6 + 20 && x < X6 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y3 + 12 && y < Y3 + 48) : 


             (array[135:132] == 4'b1000) ? (x > X6 + 20 && x < X6 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X6 + 45 && x < X6 + 52 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                         
             (array[135:132] == 4'b1001) ?  (x > X6 + 20 && x < X6 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                        (x > X6 + 20 && x < X6 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X6 + 45 && x < X6 + 52 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                        (x > X6 + 20 && x < X6 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        0;

assign num[34] = (array[139:136] == 4'b0001) ? (x > X7 + 30 && x < X7 + 42 && y > Y3 + 6 && y < Y3 + 48) :



              (array[139:136] == 4'b0010) ? ((x > X7 + 20 && x < X7 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y3 + 30 && y < Y3 + 42)) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y3 + 42 && y < Y3 + 48):


                
              (array[139:136] == 4'b0011) ? (x > X7 + 20 && x < X7 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y3 + 42 && y < Y3 + 48):

  
              (array[139:136] == 4'b0100) ? (x > X7 + 20 && x < X7 + 27 && y > Y3 + 6 && y < Y3 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y3 + 6 && y < Y3 + 48): 


             (array[139:136] == 4'b0101) ? (x > X7 + 20 && x < X7 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y3 + 42 && y < Y3 + 48) :

             (array[139:136] == 4'b0110) ? (x > X7 + 20 && x < X7 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        
             (array[139:136] == 4'b0111) ?   (x > X7 + 20 && x < X7 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y3 + 12 && y < Y3 + 48) : 


             (array[139:136] == 4'b1000) ? (x > X7 + 20 && x < X7 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X7 + 45 && x < X7 + 52 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                         
             (array[139:136] == 4'b1001) ?  (x > X7 + 20 && x < X7 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                        (x > X7 + 20 && x < X7 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X7 + 45 && x < X7 + 52 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                        (x > X7 + 20 && x < X7 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        0;

assign num[35] = (array[143:140] == 4'b0001) ? (x > X8 + 30 && x < X8 + 42 && y > Y3 + 6 && y < Y3 + 48) :



              (array[143:140] == 4'b0010) ? ((x > X8 + 20 && x < X8 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y3 + 30 && y < Y3 + 42)) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y3 + 42 && y < Y3 + 48):


                
              (array[143:140] == 4'b0011) ? (x > X8 + 20 && x < X8 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y3 + 12 && y < Y3 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y3 + 42 && y < Y3 + 48):

  
              (array[143:140] == 4'b0100) ? (x > X8 + 20 && x < X8 + 27 && y > Y3 + 6 && y < Y3 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y3 + 6 && y < Y3 + 48): 


             (array[143:140] == 4'b0101) ? (x > X8 + 20 && x < X8 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y3 + 42 && y < Y3 + 48) :

             (array[143:140] == 4'b0110) ? (x > X8 + 20 && x < X8 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y3 + 24 && y < Y3 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y3 + 30 && y < Y3 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        
             (array[143:140] == 4'b0111) ?   (x > X8 + 20 && x < X8 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y3 + 12 && y < Y3 + 48) : 


             (array[143:140] == 4'b1000) ? (x > X8 + 20 && x < X8 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X8 + 45 && x < X8 + 52 && y > Y3 + 12 && y < Y3 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                         
             (array[143:140] == 4'b1001) ?  (x > X8 + 20 && x < X8 + 52 && y > Y3 + 6 && y < Y3 + 12) || 
                                        (x > X8 + 20 && x < X8 + 27 && y > Y3 + 12 && y < Y3 + 24) || 
                                        (x > X8 + 45 && x < X8 + 52 && y > Y3 + 12 && y < Y3 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y3 + 24 && y < Y3 + 30) ||
                                        (x > X8 + 20 && x < X8 + 52 && y > Y3 + 42 && y < Y3 + 48) : 
                                        0;
                                        
                                        
                                        
  assign num[72] = (array[291:288] == 4'b0001) ? (x > X0 + 30 && x < X0 + 42 && y > Y8 + 6 && y < Y8 + 48) :



              (array[291:288] == 4'b0010) ? ((x > X0 + 20 && x < X0 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y8 + 30 && y < Y8 + 42)) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y8 + 42 && y < Y8 + 48):


                
              (array[291:288] == 4'b0011) ? (x > X0 + 20 && x < X0 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y8 + 42 && y < Y8 + 48):

  
              (array[291:288] == 4'b0100) ? (x > X0 + 20 && x < X0 + 27 && y > Y8 + 6 && y < Y8 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y8 + 6 && y < Y8 + 48): 


             (array[291:288] == 4'b0101) ? (x > X0 + 20 && x < X0 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y8 + 42 && y < Y8 + 48) :

             (array[291:288] == 4'b0110) ? (x > X0 + 20 && x < X0 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        
             (array[291:288] == 4'b0111) ?   (x > X0 + 20 && x < X0 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y8 + 12 && y < Y8 + 48) : 


             (array[291:288] == 4'b1000) ? (x > X0 + 20 && x < X0 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X0 + 45 && x < X0 + 52 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                         
             (array[291:288] == 4'b1001) ?  (x > X0 + 20 && x < X0 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                        (x > X0 + 20 && x < X0 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X0 + 45 && x < X0 + 52 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                        (x > X0 + 20 && x < X0 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        0;

assign num[73] = (array[295:292] == 4'b0001) ? (x > X1 + 30 && x < X1 + 42 && y > Y8 + 6 && y < Y8 + 48) :



              (array[295:292] == 4'b0010) ? ((x > X1 + 20 && x < X1 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y8 + 30 && y < Y8 + 42)) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y8 + 42 && y < Y8 + 48):


                
              (array[295:292] == 4'b0011) ? (x > X1 + 20 && x < X1 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y8 + 42 && y < Y8 + 48):

  
              (array[295:292] == 4'b0100) ? (x > X1 + 20 && x < X1 + 27 && y > Y8 + 6 && y < Y8 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y8 + 6 && y < Y8 + 48): 


             (array[295:292] == 4'b0101) ? (x > X1 + 20 && x < X1 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y8 + 42 && y < Y8 + 48) :

             (array[295:292] == 4'b0110) ? (x > X1 + 20 && x < X1 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        
             (array[295:292] == 4'b0111) ?   (x > X1 + 20 && x < X1 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y8 + 12 && y < Y8 + 48) : 


             (array[295:292] == 4'b1000) ? (x > X1 + 20 && x < X1 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X1 + 45 && x < X1 + 52 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                         
             (array[295:292] == 4'b1001) ?  (x > X1 + 20 && x < X1 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                        (x > X1 + 20 && x < X1 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X1 + 45 && x < X1 + 52 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                        (x > X1 + 20 && x < X1 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        0;

assign num[74] = (array[299:296] == 4'b0001) ? (x > X2 + 30 && x < X2 + 42 && y > Y8 + 6 && y < Y8 + 48) :



              (array[299:296] == 4'b0010) ? ((x > X2 + 20 && x < X2 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y8 + 30 && y < Y8 + 42)) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y8 + 42 && y < Y8 + 48):


                
              (array[299:296] == 4'b0011) ? (x > X2 + 20 && x < X2 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y8 + 42 && y < Y8 + 48):

  
              (array[299:296] == 4'b0100) ? (x > X2 + 20 && x < X2 + 27 && y > Y8 + 6 && y < Y8 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y8 + 6 && y < Y8 + 48): 


             (array[299:296] == 4'b0101) ? (x > X2 + 20 && x < X2 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y8 + 42 && y < Y8 + 48) :

             (array[299:296] == 4'b0110) ? (x > X2 + 20 && x < X2 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        
             (array[299:296] == 4'b0111) ?   (x > X2 + 20 && x < X2 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y8 + 12 && y < Y8 + 48) : 


             (array[299:296] == 4'b1000) ? (x > X2 + 20 && x < X2 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X2 + 45 && x < X2 + 52 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                         
             (array[299:296] == 4'b1001) ?  (x > X2 + 20 && x < X2 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                        (x > X2 + 20 && x < X2 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X2 + 45 && x < X2 + 52 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                        (x > X2 + 20 && x < X2 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        0;

assign num[75] = (array[303:300] == 4'b0001) ? (x > X3 + 30 && x < X3 + 42 && y > Y8 + 6 && y < Y8 + 48) :



              (array[303:300] == 4'b0010) ? ((x > X3 + 20 && x < X3 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y8 + 30 && y < Y8 + 42)) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y8 + 42 && y < Y8 + 48):


                
              (array[303:300] == 4'b0011) ? (x > X3 + 20 && x < X3 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y8 + 42 && y < Y8 + 48):

  
              (array[303:300] == 4'b0100) ? (x > X3 + 20 && x < X3 + 27 && y > Y8 + 6 && y < Y8 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y8 + 6 && y < Y8 + 48): 


             (array[303:300] == 4'b0101) ? (x > X3 + 20 && x < X3 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y8 + 42 && y < Y8 + 48) :

             (array[303:300] == 4'b0110) ? (x > X3 + 20 && x < X3 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        
             (array[303:300] == 4'b0111) ?   (x > X3 + 20 && x < X3 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y8 + 12 && y < Y8 + 48) : 


             (array[303:300] == 4'b1000) ? (x > X3 + 20 && x < X3 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X3 + 45 && x < X3 + 52 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                         
             (array[303:300] == 4'b1001) ?  (x > X3 + 20 && x < X3 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                        (x > X3 + 20 && x < X3 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X3 + 45 && x < X3 + 52 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                        (x > X3 + 20 && x < X3 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        0;

assign num[76] = (array[307:304] == 4'b0001) ? (x > X4 + 30 && x < X4 + 42 && y > Y8 + 6 && y < Y8 + 48) :



              (array[307:304] == 4'b0010) ? ((x > X4 + 20 && x < X4 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y8 + 30 && y < Y8 + 42)) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y8 + 42 && y < Y8 + 48):


                
              (array[307:304] == 4'b0011) ? (x > X4 + 20 && x < X4 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y8 + 42 && y < Y8 + 48):

  
              (array[307:304] == 4'b0100) ? (x > X4 + 20 && x < X4 + 27 && y > Y8 + 6 && y < Y8 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y8 + 6 && y < Y8 + 48): 


             (array[307:304] == 4'b0101) ? (x > X4 + 20 && x < X4 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y8 + 42 && y < Y8 + 48) :

             (array[307:304] == 4'b0110) ? (x > X4 + 20 && x < X4 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        
             (array[307:304] == 4'b0111) ?   (x > X4 + 20 && x < X4 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y8 + 12 && y < Y8 + 48) : 


             (array[307:304] == 4'b1000) ? (x > X4 + 20 && x < X4 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X4 + 45 && x < X4 + 52 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                         
             (array[307:304] == 4'b1001) ?  (x > X4 + 20 && x < X4 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                        (x > X4 + 20 && x < X4 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X4 + 45 && x < X4 + 52 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                        (x > X4 + 20 && x < X4 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        0;

assign num[77] = (array[311:308] == 4'b0001) ? (x > X5 + 30 && x < X5 + 42 && y > Y8 + 6 && y < Y8 + 48) :



              (array[311:308] == 4'b0010) ? ((x > X5 + 20 && x < X5 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y8 + 30 && y < Y8 + 42)) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y8 + 42 && y < Y8 + 48):


                
              (array[311:308] == 4'b0011) ? (x > X5 + 20 && x < X5 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y8 + 42 && y < Y8 + 48):

  
              (array[311:308] == 4'b0100) ? (x > X5 + 20 && x < X5 + 27 && y > Y8 + 6 && y < Y8 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y8 + 6 && y < Y8 + 48): 


             (array[311:308] == 4'b0101) ? (x > X5 + 20 && x < X5 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y8 + 42 && y < Y8 + 48) :

             (array[311:308] == 4'b0110) ? (x > X5 + 20 && x < X5 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        
             (array[311:308] == 4'b0111) ?   (x > X5 + 20 && x < X5 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y8 + 12 && y < Y8 + 48) : 


             (array[311:308] == 4'b1000) ? (x > X5 + 20 && x < X5 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X5 + 45 && x < X5 + 52 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                         
             (array[311:308] == 4'b1001) ?  (x > X5 + 20 && x < X5 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                        (x > X5 + 20 && x < X5 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X5 + 45 && x < X5 + 52 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                        (x > X5 + 20 && x < X5 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        0;

assign num[78] = (array[315:312] == 4'b0001) ? (x > X6 + 30 && x < X6 + 42 && y > Y8 + 6 && y < Y8 + 48) :



              (array[315:312] == 4'b0010) ? ((x > X6 + 20 && x < X6 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y8 + 30 && y < Y8 + 42)) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y8 + 42 && y < Y8 + 48):


                
              (array[315:312] == 4'b0011) ? (x > X6 + 20 && x < X6 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y8 + 42 && y < Y8 + 48):

  
              (array[315:312] == 4'b0100) ? (x > X6 + 20 && x < X6 + 27 && y > Y8 + 6 && y < Y8 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y8 + 6 && y < Y8 + 48): 


             (array[315:312] == 4'b0101) ? (x > X6 + 20 && x < X6 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y8 + 42 && y < Y8 + 48) :

             (array[315:312] == 4'b0110) ? (x > X6 + 20 && x < X6 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        
             (array[315:312] == 4'b0111) ?   (x > X6 + 20 && x < X6 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y8 + 12 && y < Y8 + 48) : 


             (array[315:312] == 4'b1000) ? (x > X6 + 20 && x < X6 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X6 + 45 && x < X6 + 52 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                         
             (array[315:312] == 4'b1001) ?  (x > X6 + 20 && x < X6 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                        (x > X6 + 20 && x < X6 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X6 + 45 && x < X6 + 52 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                        (x > X6 + 20 && x < X6 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        0;

assign num[79] = (array[319:316] == 4'b0001) ? (x > X7 + 30 && x < X7 + 42 && y > Y8 + 6 && y < Y8 + 48) :



              (array[319:316] == 4'b0010) ? ((x > X7 + 20 && x < X7 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y8 + 30 && y < Y8 + 42)) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y8 + 42 && y < Y8 + 48):


                
              (array[319:316] == 4'b0011) ? (x > X7 + 20 && x < X7 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y8 + 42 && y < Y8 + 48):

  
              (array[319:316] == 4'b0100) ? (x > X7 + 20 && x < X7 + 27 && y > Y8 + 6 && y < Y8 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y8 + 6 && y < Y8 + 48): 


             (array[319:316] == 4'b0101) ? (x > X7 + 20 && x < X7 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y8 + 42 && y < Y8 + 48) :

             (array[319:316] == 4'b0110) ? (x > X7 + 20 && x < X7 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        
             (array[319:316] == 4'b0111) ?   (x > X7 + 20 && x < X7 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y8 + 12 && y < Y8 + 48) : 


             (array[319:316] == 4'b1000) ? (x > X7 + 20 && x < X7 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X7 + 45 && x < X7 + 52 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                         
             (array[319:316] == 4'b1001) ?  (x > X7 + 20 && x < X7 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                        (x > X7 + 20 && x < X7 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X7 + 45 && x < X7 + 52 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                        (x > X7 + 20 && x < X7 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        0;

assign num[80] = (array[323:320] == 4'b0001) ? (x > X8 + 30 && x < X8 + 42 && y > Y8 + 6 && y < Y8 + 48) :



              (array[323:320] == 4'b0010) ? ((x > X8 + 20 && x < X8 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y8 + 30 && y < Y8 + 42)) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y8 + 42 && y < Y8 + 48):


                
              (array[323:320] == 4'b0011) ? (x > X8 + 20 && x < X8 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y8 + 12 && y < Y8 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y8 + 42 && y < Y8 + 48):

  
              (array[323:320] == 4'b0100) ? (x > X8 + 20 && x < X8 + 27 && y > Y8 + 6 && y < Y8 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y8 + 6 && y < Y8 + 48): 


             (array[323:320] == 4'b0101) ? (x > X8 + 20 && x < X8 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y8 + 42 && y < Y8 + 48) :

             (array[323:320] == 4'b0110) ? (x > X8 + 20 && x < X8 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y8 + 24 && y < Y8 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y8 + 30 && y < Y8 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        
             (array[323:320] == 4'b0111) ?   (x > X8 + 20 && x < X8 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y8 + 12 && y < Y8 + 48) : 


             (array[323:320] == 4'b1000) ? (x > X8 + 20 && x < X8 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X8 + 45 && x < X8 + 52 && y > Y8 + 12 && y < Y8 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                         
             (array[323:320] == 4'b1001) ?  (x > X8 + 20 && x < X8 + 52 && y > Y8 + 6 && y < Y8 + 12) || 
                                        (x > X8 + 20 && x < X8 + 27 && y > Y8 + 12 && y < Y8 + 24) || 
                                        (x > X8 + 45 && x < X8 + 52 && y > Y8 + 12 && y < Y8 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y8 + 24 && y < Y8 + 30) ||
                                        (x > X8 + 20 && x < X8 + 52 && y > Y8 + 42 && y < Y8 + 48) : 
                                        0;
                                        
                                        
                                        
                                        
                                                assign num[45] = (array[183:180] == 4'b0001) ? (x > X0 + 30 && x < X0 + 42 && y > Y5 + 6 && y < Y5 + 48) :



              (array[183:180] == 4'b0010) ? ((x > X0 + 20 && x < X0 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y5 + 30 && y < Y5 + 42)) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y5 + 42 && y < Y5 + 48):

                
              (array[183:180] == 4'b0011) ? (x > X0 + 20 && x < X0 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y5 + 42 && y < Y5 + 48):

  
              (array[183:180] == 4'b0100) ? (x > X0 + 20 && x < X0 + 27 && y > Y5 + 6 && y < Y5 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y5 + 6 && y < Y5 + 48): 


             (array[183:180] == 4'b0101) ? (x > X0 + 20 && x < X0 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y5 + 42 && y < Y5 + 48) :

             (array[183:180] == 4'b0110) ? (x > X0 + 20 && x < X0 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        
             (array[183:180] == 4'b0111) ?   (x > X0 + 20 && x < X0 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y5 + 12 && y < Y5 + 48) : 


             (array[183:180] == 4'b1000) ? (x > X0 + 20 && x < X0 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X0 + 45 && x < X0 + 52 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                         
             (array[183:180] == 4'b1001) ?  (x > X0 + 20 && x < X0 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                        (x > X0 + 20 && x < X0 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X0 + 45 && x < X0 + 52 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                        (x > X0 + 20 && x < X0 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        0;      
                
  
        assign num[46] = (array[187:184] == 4'b0001) ? (x > X1 + 30 && x < X1 + 42 && y > Y5 + 6 && y < Y5 + 48) :



              (array[187:184] == 4'b0010) ? ((x > X1 + 20 && x < X1 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y5 + 30 && y < Y5 + 42)) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y5 + 42 && y < Y5 + 48):

                
              (array[187:184] == 4'b0011) ? (x > X1 + 20 && x < X1 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y5 + 42 && y < Y5 + 48):

  
              (array[187:184] == 4'b0100) ? (x > X1 + 20 && x < X1 + 27 && y > Y5 + 6 && y < Y5 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y5 + 6 && y < Y5 + 48): 


             (array[187:184] == 4'b0101) ? (x > X1 + 20 && x < X1 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y5 + 42 && y < Y5 + 48) :

             (array[187:184] == 4'b0110) ? (x > X1 + 20 && x < X1 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        
             (array[187:184] == 4'b0111) ?   (x > X1 + 20 && x < X1 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y5 + 12 && y < Y5 + 48) : 


             (array[187:184] == 4'b1000) ? (x > X1 + 20 && x < X1 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X1 + 45 && x < X1 + 52 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                         
             (array[187:184] == 4'b1001) ?  (x > X1 + 20 && x < X1 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                        (x > X1 + 20 && x < X1 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X1 + 45 && x < X1 + 52 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                        (x > X1 + 20 && x < X1 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        0;      
                

        assign num[47] = (array[191:188] == 4'b0001) ? (x > X2 + 30 && x < X2 + 42 && y > Y5 + 6 && y < Y5 + 48) :



              (array[191:188] == 4'b0010) ? ((x > X2 + 20 && x < X2 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y5 + 30 && y < Y5 + 42)) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y5 + 42 && y < Y5 + 48):

                
              (array[191:188] == 4'b0011) ? (x > X2 + 20 && x < X2 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y5 + 42 && y < Y5 + 48):

  
              (array[191:188] == 4'b0100) ? (x > X2 + 20 && x < X2 + 27 && y > Y5 + 6 && y < Y5 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y5 + 6 && y < Y5 + 48): 


             (array[191:188] == 4'b0101) ? (x > X2 + 20 && x < X2 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y5 + 42 && y < Y5 + 48) :

             (array[191:188] == 4'b0110) ? (x > X2 + 20 && x < X2 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        
             (array[191:188] == 4'b0111) ?   (x > X2 + 20 && x < X2 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y5 + 12 && y < Y5 + 48) : 


             (array[191:188] == 4'b1000) ? (x > X2 + 20 && x < X2 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X2 + 45 && x < X2 + 52 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                         
             (array[191:188] == 4'b1001) ?  (x > X2 + 20 && x < X2 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                        (x > X2 + 20 && x < X2 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X2 + 45 && x < X2 + 52 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                        (x > X2 + 20 && x < X2 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        0;

        assign num[48] = (array[195:192] == 4'b0001) ? (x > X3 + 30 && x < X3 + 42 && y > Y5 + 6 && y < Y5 + 48) :



              (array[195:192] == 4'b0010) ? ((x > X3 + 20 && x < X3 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y5 + 30 && y < Y5 + 42)) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y5 + 42 && y < Y5 + 48):

                
              (array[195:192] == 4'b0011) ? (x > X3 + 20 && x < X3 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y5 + 42 && y < Y5 + 48):

  
              (array[195:192] == 4'b0100) ? (x > X3 + 20 && x < X3 + 27 && y > Y5 + 6 && y < Y5 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y5 + 6 && y < Y5 + 48): 


             (array[195:192] == 4'b0101) ? (x > X3 + 20 && x < X3 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y5 + 42 && y < Y5 + 48) :

             (array[195:192] == 4'b0110) ? (x > X3 + 20 && x < X3 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        
             (array[195:192] == 4'b0111) ?   (x > X3 + 20 && x < X3 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y5 + 12 && y < Y5 + 48) : 


             (array[195:192] == 4'b1000) ? (x > X3 + 20 && x < X3 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X3 + 45 && x < X3 + 52 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                         
             (array[195:192] == 4'b1001) ?  (x > X3 + 20 && x < X3 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                        (x > X3 + 20 && x < X3 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X3 + 45 && x < X3 + 52 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                        (x > X3 + 20 && x < X3 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        0;

        assign num[49] = (array[199:196] == 4'b0001) ? (x > X4 + 30 && x < X4 + 42 && y > Y5 + 6 && y < Y5 + 48) :



              (array[199:196] == 4'b0010) ? ((x > X4 + 20 && x < X4 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y5 + 30 && y < Y5 + 42)) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y5 + 42 && y < Y5 + 48):

                
              (array[199:196] == 4'b0011) ? (x > X4 + 20 && x < X4 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y5 + 42 && y < Y5 + 48):

  
              (array[199:196] == 4'b0100) ? (x > X4 + 20 && x < X4 + 27 && y > Y5 + 6 && y < Y5 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y5 + 6 && y < Y5 + 48): 


             (array[199:196] == 4'b0101) ? (x > X4 + 20 && x < X4 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y5 + 42 && y < Y5 + 48) :

             (array[199:196] == 4'b0110) ? (x > X4 + 20 && x < X4 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        
             (array[199:196] == 4'b0111) ?   (x > X4 + 20 && x < X4 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y5 + 12 && y < Y5 + 48) : 


             (array[199:196] == 4'b1000) ? (x > X4 + 20 && x < X4 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X4 + 45 && x < X4 + 52 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                         
             (array[199:196] == 4'b1001) ?  (x > X4 + 20 && x < X4 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                        (x > X4 + 20 && x < X4 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X4 + 45 && x < X4 + 52 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                        (x > X4 + 20 && x < X4 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        0;



        assign num[50] = (array[203:200] == 4'b0001) ? (x > X5 + 30 && x < X5 + 42 && y > Y5 + 6 && y < Y5 + 48) :



              (array[203:200] == 4'b0010) ? ((x > X5 + 20 && x < X5 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y5 + 30 && y < Y5 + 42)) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y5 + 42 && y < Y5 + 48):

                
              (array[203:200] == 4'b0011) ? (x > X5 + 20 && x < X5 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y5 + 42 && y < Y5 + 48):

  
              (array[203:200] == 4'b0100) ? (x > X5 + 20 && x < X5 + 27 && y > Y5 + 6 && y < Y5 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y5 + 6 && y < Y5 + 48): 


             (array[203:200] == 4'b0101) ? (x > X5 + 20 && x < X5 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y5 + 42 && y < Y5 + 48) :

             (array[203:200] == 4'b0110) ? (x > X5 + 20 && x < X5 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        
             (array[203:200] == 4'b0111) ?   (x > X5 + 20 && x < X5 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y5 + 12 && y < Y5 + 48) : 


             (array[203:200] == 4'b1000) ? (x > X5 + 20 && x < X5 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X5 + 45 && x < X5 + 52 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                         
             (array[203:200] == 4'b1001) ?  (x > X5 + 20 && x < X5 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                        (x > X5 + 20 && x < X5 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X5 + 45 && x < X5 + 52 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                        (x > X5 + 20 && x < X5 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        0;


        assign num[51] = (array[207:204] == 4'b0001) ? (x > X6 + 30 && x < X6 + 42 && y > Y5 + 6 && y < Y5 + 48) :



              (array[207:204] == 4'b0010) ? ((x > X6 + 20 && x < X6 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y5 + 30 && y < Y5 + 42)) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y5 + 42 && y < Y5 + 48):

                
              (array[207:204] == 4'b0011) ? (x > X6 + 20 && x < X6 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y5 + 42 && y < Y5 + 48):

  
              (array[207:204] == 4'b0100) ? (x > X6 + 20 && x < X6 + 27 && y > Y5 + 6 && y < Y5 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y5 + 6 && y < Y5 + 48): 


             (array[207:204] == 4'b0101) ? (x > X6 + 20 && x < X6 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y5 + 42 && y < Y5 + 48) :

             (array[207:204] == 4'b0110) ? (x > X6 + 20 && x < X6 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        
             (array[207:204] == 4'b0111) ?   (x > X6 + 20 && x < X6 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y5 + 12 && y < Y5 + 48) : 


             (array[207:204] == 4'b1000) ? (x > X6 + 20 && x < X6 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X6 + 45 && x < X6 + 52 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                         
             (array[207:204] == 4'b1001) ?  (x > X6 + 20 && x < X6 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                        (x > X6 + 20 && x < X6 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X6 + 45 && x < X6 + 52 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                        (x > X6 + 20 && x < X6 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        0;

        assign num[52] = (array[211:208] == 4'b0001) ? (x > X7 + 30 && x < X7 + 42 && y > Y5 + 6 && y < Y5 + 48) :



              (array[211:208] == 4'b0010) ? ((x > X7 + 20 && x < X7 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y5 + 30 && y < Y5 + 42)) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y5 + 42 && y < Y5 + 48):

                
              (array[211:208] == 4'b0011) ? (x > X7 + 20 && x < X7 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y5 + 42 && y < Y5 + 48):

  
              (array[211:208] == 4'b0100) ? (x > X7 + 20 && x < X7 + 27 && y > Y5 + 6 && y < Y5 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y5 + 6 && y < Y5 + 48): 


             (array[211:208] == 4'b0101) ? (x > X7 + 20 && x < X7 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y5 + 42 && y < Y5 + 48) :

             (array[211:208] == 4'b0110) ? (x > X7 + 20 && x < X7 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        
             (array[211:208] == 4'b0111) ?   (x > X7 + 20 && x < X7 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y5 + 12 && y < Y5 + 48) : 


             (array[211:208] == 4'b1000) ? (x > X7 + 20 && x < X7 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X7 + 45 && x < X7 + 52 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                         
             (array[211:208] == 4'b1001) ?  (x > X7 + 20 && x < X7 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                        (x > X7 + 20 && x < X7 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X7 + 45 && x < X7 + 52 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                        (x > X7 + 20 && x < X7 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        0;



        assign num[53] = (array[215:212] == 4'b0001) ? (x > X8 + 30 && x < X8 + 42 && y > Y5 + 6 && y < Y5 + 48) :



              (array[215:212] == 4'b0010) ? ((x > X8 + 20 && x < X8 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y5 + 30 && y < Y5 + 42)) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y5 + 42 && y < Y5 + 48):

                
              (array[215:212] == 4'b0011) ? (x > X8 + 20 && x < X8 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y5 + 12 && y < Y5 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y5 + 42 && y < Y5 + 48):

  
              (array[215:212] == 4'b0100) ? (x > X8 + 20 && x < X8 + 27 && y > Y5 + 6 && y < Y5 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y5 + 6 && y < Y5 + 48): 


             (array[215:212] == 4'b0101) ? (x > X8 + 20 && x < X8 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y5 + 42 && y < Y5 + 48) :

             (array[215:212] == 4'b0110) ? (x > X8 + 20 && x < X8 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y5 + 24 && y < Y5 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y5 + 30 && y < Y5 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        
             (array[215:212] == 4'b0111) ?   (x > X8 + 20 && x < X8 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y5 + 12 && y < Y5 + 48) : 


             (array[215:212] == 4'b1000) ? (x > X8 + 20 && x < X8 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X8 + 45 && x < X8 + 52 && y > Y5 + 12 && y < Y5 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                         
             (array[215:212] == 4'b1001) ?  (x > X8 + 20 && x < X8 + 52 && y > Y5 + 6 && y < Y5 + 12) || 
                                        (x > X8 + 20 && x < X8 + 27 && y > Y5 + 12 && y < Y5 + 24) || 
                                        (x > X8 + 45 && x < X8 + 52 && y > Y5 + 12 && y < Y5 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y5 + 24 && y < Y5 + 30) ||
                                        (x > X8 + 20 && x < X8 + 52 && y > Y5 + 42 && y < Y5 + 48) : 
                                        0;
                                        
                                        
                                        assign num[36] = (array[147:144] == 4'b0001) ? (x > X0 + 30 && x < X0 + 42 && y > Y4 + 6 && y < Y4 + 48) :



              (array[147:144] == 4'b0010) ? ((x > X0 + 20 && x < X0 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y4 + 30 && y < Y4 + 42)) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y4 + 42 && y < Y4 + 48):


                
              (array[147:144] == 4'b0011) ? (x > X0 + 20 && x < X0 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y4 + 42 && y < Y4 + 48):

  
              (array[147:144] == 4'b0100) ? (x > X0 + 20 && x < X0 + 27 && y > Y4 + 6 && y < Y4 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y4 + 6 && y < Y4 + 48): 


             (array[147:144] == 4'b0101) ? (x > X0 + 20 && x < X0 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y4 + 42 && y < Y4 + 48) :

             (array[147:144] == 4'b0110) ? (x > X0 + 20 && x < X0 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        
             (array[147:144] == 4'b0111) ?   (x > X0 + 20 && x < X0 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y4 + 12 && y < Y4 + 48) : 


             (array[147:144] == 4'b1000) ? (x > X0 + 20 && x < X0 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X0 + 45 && x < X0 + 52 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                         
             (array[147:144] == 4'b1001) ?  (x > X0 + 20 && x < X0 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                        (x > X0 + 20 && x < X0 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X0 + 45 && x < X0 + 52 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                        (x > X0 + 20 && x < X0 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        0;

assign num[37] = (array[151:148] == 4'b0001) ? (x > X1 + 30 && x < X1 + 42 && y > Y4 + 6 && y < Y4 + 48) :



              (array[151:148] == 4'b0010) ? ((x > X1 + 20 && x < X1 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y4 + 30 && y < Y4 + 42)) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y4 + 42 && y < Y4 + 48):


                
              (array[151:148] == 4'b0011) ? (x > X1 + 20 && x < X1 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y4 + 42 && y < Y4 + 48):

  
              (array[151:148] == 4'b0100) ? (x > X1 + 20 && x < X1 + 27 && y > Y4 + 6 && y < Y4 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y4 + 6 && y < Y4 + 48): 


             (array[151:148] == 4'b0101) ? (x > X1 + 20 && x < X1 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y4 + 42 && y < Y4 + 48) :

             (array[151:148] == 4'b0110) ? (x > X1 + 20 && x < X1 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        
             (array[151:148] == 4'b0111) ?   (x > X1 + 20 && x < X1 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y4 + 12 && y < Y4 + 48) : 


             (array[151:148] == 4'b1000) ? (x > X1 + 20 && x < X1 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X1 + 45 && x < X1 + 52 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                         
             (array[151:148] == 4'b1001) ?  (x > X1 + 20 && x < X1 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                        (x > X1 + 20 && x < X1 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X1 + 45 && x < X1 + 52 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                        (x > X1 + 20 && x < X1 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        0;

assign num[38] = (array[155:152] == 4'b0001) ? (x > X2 + 30 && x < X2 + 42 && y > Y4 + 6 && y < Y4 + 48) :



              (array[155:152] == 4'b0010) ? ((x > X2 + 20 && x < X2 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y4 + 30 && y < Y4 + 42)) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y4 + 42 && y < Y4 + 48):


                
              (array[155:152] == 4'b0011) ? (x > X2 + 20 && x < X2 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y4 + 42 && y < Y4 + 48):

  
              (array[155:152] == 4'b0100) ? (x > X2 + 20 && x < X2 + 27 && y > Y4 + 6 && y < Y4 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y4 + 6 && y < Y4 + 48): 


             (array[155:152] == 4'b0101) ? (x > X2 + 20 && x < X2 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y4 + 42 && y < Y4 + 48) :

             (array[155:152] == 4'b0110) ? (x > X2 + 20 && x < X2 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        
             (array[155:152] == 4'b0111) ?   (x > X2 + 20 && x < X2 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y4 + 12 && y < Y4 + 48) : 


             (array[155:152] == 4'b1000) ? (x > X2 + 20 && x < X2 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X2 + 45 && x < X2 + 52 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                         
             (array[155:152] == 4'b1001) ?  (x > X2 + 20 && x < X2 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                        (x > X2 + 20 && x < X2 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X2 + 45 && x < X2 + 52 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                        (x > X2 + 20 && x < X2 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        0;
assign num[39] = (array[159:156] == 4'b0001) ? (x > X3 + 30 && x < X3 + 42 && y > Y4 + 6 && y < Y4 + 48) :



              (array[159:156] == 4'b0010) ? ((x > X3 + 20 && x < X3 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y4 + 30 && y < Y4 + 42)) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y4 + 42 && y < Y4 + 48):


                
              (array[159:156] == 4'b0011) ? (x > X3 + 20 && x < X3 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y4 + 42 && y < Y4 + 48):

  
              (array[159:156] == 4'b0100) ? (x > X3 + 20 && x < X3 + 27 && y > Y4 + 6 && y < Y4 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y4 + 6 && y < Y4 + 48): 


             (array[159:156] == 4'b0101) ? (x > X3 + 20 && x < X3 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y4 + 42 && y < Y4 + 48) :

             (array[159:156] == 4'b0110) ? (x > X3 + 20 && x < X3 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        
             (array[159:156] == 4'b0111) ?   (x > X3 + 20 && x < X3 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y4 + 12 && y < Y4 + 48) : 


             (array[159:156] == 4'b1000) ? (x > X3 + 20 && x < X3 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X3 + 45 && x < X3 + 52 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                         
             (array[159:156] == 4'b1001) ?  (x > X3 + 20 && x < X3 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                        (x > X3 + 20 && x < X3 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X3 + 45 && x < X3 + 52 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                        (x > X3 + 20 && x < X3 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        0;

assign num[40] = (array[163:160] == 4'b0001) ? (x > X4 + 30 && x < X4 + 42 && y > Y4 + 6 && y < Y4 + 48) :



              (array[163:160] == 4'b0010) ? ((x > X4 + 20 && x < X4 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y4 + 30 && y < Y4 + 42)) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y4 + 42 && y < Y4 + 48):


                
              (array[163:160] == 4'b0011) ? (x > X4 + 20 && x < X4 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y4 + 42 && y < Y4 + 48):

  
              (array[163:160] == 4'b0100) ? (x > X4 + 20 && x < X4 + 27 && y > Y4 + 6 && y < Y4 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y4 + 6 && y < Y4 + 48): 


             (array[163:160] == 4'b0101) ? (x > X4 + 20 && x < X4 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y4 + 42 && y < Y4 + 48) :

             (array[163:160] == 4'b0110) ? (x > X4 + 20 && x < X4 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        
             (array[163:160] == 4'b0111) ?   (x > X4 + 20 && x < X4 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y4 + 12 && y < Y4 + 48) : 


             (array[163:160] == 4'b1000) ? (x > X4 + 20 && x < X4 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X4 + 45 && x < X4 + 52 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                         
             (array[163:160] == 4'b1001) ?  (x > X4 + 20 && x < X4 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                        (x > X4 + 20 && x < X4 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X4 + 45 && x < X4 + 52 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                        (x > X4 + 20 && x < X4 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        0;

assign num[41] = (array[167:164] == 4'b0001) ? (x > X5 + 30 && x < X5 + 42 && y > Y4 + 6 && y < Y4 + 48) :



              (array[167:164] == 4'b0010) ? ((x > X5 + 20 && x < X5 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y4 + 30 && y < Y4 + 42)) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y4 + 42 && y < Y4 + 48):


                
              (array[167:164] == 4'b0011) ? (x > X5 + 20 && x < X5 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y4 + 42 && y < Y4 + 48):

  
              (array[167:164] == 4'b0100) ? (x > X5 + 20 && x < X5 + 27 && y > Y4 + 6 && y < Y4 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y4 + 6 && y < Y4 + 48): 


             (array[167:164] == 4'b0101) ? (x > X5 + 20 && x < X5 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y4 + 42 && y < Y4 + 48) :

             (array[167:164] == 4'b0110) ? (x > X5 + 20 && x < X5 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        
             (array[167:164] == 4'b0111) ?   (x > X5 + 20 && x < X5 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y4 + 12 && y < Y4 + 48) : 


             (array[167:164] == 4'b1000) ? (x > X5 + 20 && x < X5 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X5 + 45 && x < X5 + 52 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                         
             (array[167:164] == 4'b1001) ?  (x > X5 + 20 && x < X5 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                        (x > X5 + 20 && x < X5 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X5 + 45 && x < X5 + 52 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                        (x > X5 + 20 && x < X5 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        0;

assign num[42] = (array[171:168] == 4'b0001) ? (x > X6 + 30 && x < X6 + 42 && y > Y4 + 6 && y < Y4 + 48) :



              (array[171:168] == 4'b0010) ? ((x > X6 + 20 && x < X6 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y4 + 30 && y < Y4 + 42)) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y4 + 42 && y < Y4 + 48):


                
              (array[171:168] == 4'b0011) ? (x > X6 + 20 && x < X6 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y4 + 42 && y < Y4 + 48):

  
              (array[171:168] == 4'b0100) ? (x > X6 + 20 && x < X6 + 27 && y > Y4 + 6 && y < Y4 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y4 + 6 && y < Y4 + 48): 


             (array[171:168] == 4'b0101) ? (x > X6 + 20 && x < X6 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y4 + 42 && y < Y4 + 48) :

             (array[171:168] == 4'b0110) ? (x > X6 + 20 && x < X6 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        
             (array[171:168] == 4'b0111) ?   (x > X6 + 20 && x < X6 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y4 + 12 && y < Y4 + 48) : 


             (array[171:168] == 4'b1000) ? (x > X6 + 20 && x < X6 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X6 + 45 && x < X6 + 52 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                         
             (array[171:168] == 4'b1001) ?  (x > X6 + 20 && x < X6 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                        (x > X6 + 20 && x < X6 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X6 + 45 && x < X6 + 52 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                        (x > X6 + 20 && x < X6 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        0;

assign num[43] = (array[175:172] == 4'b0001) ? (x > X7 + 30 && x < X7 + 42 && y > Y4 + 6 && y < Y4 + 48) :



              (array[175:172] == 4'b0010) ? ((x > X7 + 20 && x < X7 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y4 + 30 && y < Y4 + 42)) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y4 + 42 && y < Y4 + 48):


                
              (array[175:172] == 4'b0011) ? (x > X7 + 20 && x < X7 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y4 + 42 && y < Y4 + 48):

  
              (array[175:172] == 4'b0100) ? (x > X7 + 20 && x < X7 + 27 && y > Y4 + 6 && y < Y4 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y4 + 6 && y < Y4 + 48): 


             (array[175:172] == 4'b0101) ? (x > X7 + 20 && x < X7 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y4 + 42 && y < Y4 + 48) :

             (array[175:172] == 4'b0110) ? (x > X7 + 20 && x < X7 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        
             (array[175:172] == 4'b0111) ?   (x > X7 + 20 && x < X7 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y4 + 12 && y < Y4 + 48) : 


             (array[175:172] == 4'b1000) ? (x > X7 + 20 && x < X7 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X7 + 45 && x < X7 + 52 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                         
             (array[175:172] == 4'b1001) ?  (x > X7 + 20 && x < X7 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                        (x > X7 + 20 && x < X7 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X7 + 45 && x < X7 + 52 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                        (x > X7 + 20 && x < X7 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        0;
assign num[44] = (array[179:176] == 4'b0001) ? (x > X8 + 30 && x < X8 + 42 && y > Y4 + 6 && y < Y4 + 48) :



              (array[179:176] == 4'b0010) ? ((x > X8 + 20 && x < X8 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y4 + 30 && y < Y4 + 42)) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y4 + 42 && y < Y4 + 48):


                
              (array[179:176] == 4'b0011) ? (x > X8 + 20 && x < X8 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y4 + 12 && y < Y4 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y4 + 42 && y < Y4 + 48):

  
              (array[179:176] == 4'b0100) ? (x > X8 + 20 && x < X8 + 27 && y > Y4 + 6 && y < Y4 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y4 + 6 && y < Y4 + 48): 


             (array[179:176] == 4'b0101) ? (x > X8 + 20 && x < X8 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y4 + 42 && y < Y4 + 48) :

             (array[179:176] == 4'b0110) ? (x > X8 + 20 && x < X8 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y4 + 24 && y < Y4 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y4 + 30 && y < Y4 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        
             (array[179:176] == 4'b0111) ?   (x > X8 + 20 && x < X8 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y4 + 12 && y < Y4 + 48) : 


             (array[179:176] == 4'b1000) ? (x > X8 + 20 && x < X8 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X8 + 45 && x < X8 + 52 && y > Y4 + 12 && y < Y4 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                         
             (array[179:176] == 4'b1001) ?  (x > X8 + 20 && x < X8 + 52 && y > Y4 + 6 && y < Y4 + 12) || 
                                        (x > X8 + 20 && x < X8 + 27 && y > Y4 + 12 && y < Y4 + 24) || 
                                        (x > X8 + 45 && x < X8 + 52 && y > Y4 + 12 && y < Y4 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y4 + 24 && y < Y4 + 30) ||
                                        (x > X8 + 20 && x < X8 + 52 && y > Y4 + 42 && y < Y4 + 48) : 
                                        0;

assign num[54] = (array[219:216] == 4'b0001) ? (x > X0 + 30 && x < X0 + 42 && y > Y6 + 6 && y < Y6 + 48) :



              (array[219:216] == 4'b0010) ? ((x > X0 + 20 && x < X0 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y6 + 30 && y < Y6 + 42)) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y6 + 42 && y < Y6 + 48):


                
              (array[219:216] == 4'b0011) ? (x > X0 + 20 && x < X0 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y6 + 42 && y < Y6 + 48):

  
              (array[219:216] == 4'b0100) ? (x > X0 + 20 && x < X0 + 27 && y > Y6 + 6 && y < Y6 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y6 + 6 && y < Y6 + 48): 


             (array[219:216] == 4'b0101) ? (x > X0 + 20 && x < X0 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y6 + 42 && y < Y6 + 48) :

             (array[219:216] == 4'b0110) ? (x > X0 + 20 && x < X0 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        
             (array[219:216] == 4'b0111) ?   (x > X0 + 20 && x < X0 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y6 + 12 && y < Y6 + 48) : 


             (array[219:216] == 4'b1000) ? (x > X0 + 20 && x < X0 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X0 + 45 && x < X0 + 52 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                         
             (array[219:216] == 4'b1001) ?  (x > X0 + 20 && x < X0 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                        (x > X0 + 20 && x < X0 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X0 + 45 && x < X0 + 52 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                        (x > X0 + 20 && x < X0 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        0;

assign num[55] = (array[223:220] == 4'b0001) ? (x > X1 + 30 && x < X1 + 42 && y > Y6 + 6 && y < Y6 + 48) :



              (array[223:220] == 4'b0010) ? ((x > X1 + 20 && x < X1 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y6 + 30 && y < Y6 + 42)) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y6 + 42 && y < Y6 + 48):


                
              (array[223:220] == 4'b0011) ? (x > X1 + 20 && x < X1 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y6 + 42 && y < Y6 + 48):

  
              (array[223:220] == 4'b0100) ? (x > X1 + 20 && x < X1 + 27 && y > Y6 + 6 && y < Y6 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y6 + 6 && y < Y6 + 48): 


             (array[223:220] == 4'b0101) ? (x > X1 + 20 && x < X1 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y6 + 42 && y < Y6 + 48) :

             (array[223:220] == 4'b0110) ? (x > X1 + 20 && x < X1 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        
             (array[223:220] == 4'b0111) ?   (x > X1 + 20 && x < X1 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y6 + 12 && y < Y6 + 48) : 


             (array[223:220] == 4'b1000) ? (x > X1 + 20 && x < X1 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X1 + 45 && x < X1 + 52 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                         
             (array[223:220] == 4'b1001) ?  (x > X1 + 20 && x < X1 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                        (x > X1 + 20 && x < X1 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X1 + 45 && x < X1 + 52 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                        (x > X1 + 20 && x < X1 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        0;

assign num[56] = (array[227:224] == 4'b0001) ? (x > X2 + 30 && x < X2 + 42 && y > Y6 + 6 && y < Y6 + 48) :



              (array[227:224] == 4'b0010) ? ((x > X2 + 20 && x < X2 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y6 + 30 && y < Y6 + 42)) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y6 + 42 && y < Y6 + 48):


                
              (array[227:224] == 4'b0011) ? (x > X2 + 20 && x < X2 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y6 + 42 && y < Y6 + 48):

  
              (array[227:224] == 4'b0100) ? (x > X2 + 20 && x < X2 + 27 && y > Y6 + 6 && y < Y6 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y6 + 6 && y < Y6 + 48): 


             (array[227:224] == 4'b0101) ? (x > X2 + 20 && x < X2 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y6 + 42 && y < Y6 + 48) :

             (array[227:224] == 4'b0110) ? (x > X2 + 20 && x < X2 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        
             (array[227:224] == 4'b0111) ?   (x > X2 + 20 && x < X2 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y6 + 12 && y < Y6 + 48) : 


             (array[227:224] == 4'b1000) ? (x > X2 + 20 && x < X2 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X2 + 45 && x < X2 + 52 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                         
             (array[227:224] == 4'b1001) ?  (x > X2 + 20 && x < X2 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                        (x > X2 + 20 && x < X2 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X2 + 45 && x < X2 + 52 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                        (x > X2 + 20 && x < X2 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        0;

assign num[57] = (array[231:228] == 4'b0001) ? (x > X3 + 30 && x < X3 + 42 && y > Y6 + 6 && y < Y6 + 48) :



              (array[231:228] == 4'b0010) ? ((x > X3 + 20 && x < X3 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y6 + 30 && y < Y6 + 42)) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y6 + 42 && y < Y6 + 48):


                
              (array[231:228] == 4'b0011) ? (x > X3 + 20 && x < X3 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y6 + 42 && y < Y6 + 48):

  
              (array[231:228] == 4'b0100) ? (x > X3 + 20 && x < X3 + 27 && y > Y6 + 6 && y < Y6 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y6 + 6 && y < Y6 + 48): 


             (array[231:228] == 4'b0101) ? (x > X3 + 20 && x < X3 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y6 + 42 && y < Y6 + 48) :

             (array[231:228] == 4'b0110) ? (x > X3 + 20 && x < X3 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        
             (array[231:228] == 4'b0111) ?   (x > X3 + 20 && x < X3 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y6 + 12 && y < Y6 + 48) : 


             (array[231:228] == 4'b1000) ? (x > X3 + 20 && x < X3 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X3 + 45 && x < X3 + 52 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                         
             (array[231:228] == 4'b1001) ?  (x > X3 + 20 && x < X3 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                        (x > X3 + 20 && x < X3 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X3 + 45 && x < X3 + 52 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                        (x > X3 + 20 && x < X3 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        0;

assign num[58] = (array[235:232] == 4'b0001) ? (x > X4 + 30 && x < X4 + 42 && y > Y6 + 6 && y < Y6 + 48) :



              (array[235:232] == 4'b0010) ? ((x > X4 + 20 && x < X4 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y6 + 30 && y < Y6 + 42)) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y6 + 42 && y < Y6 + 48):


                
              (array[235:232] == 4'b0011) ? (x > X4 + 20 && x < X4 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y6 + 42 && y < Y6 + 48):

  
              (array[235:232] == 4'b0100) ? (x > X4 + 20 && x < X4 + 27 && y > Y6 + 6 && y < Y6 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y6 + 6 && y < Y6 + 48): 


             (array[235:232] == 4'b0101) ? (x > X4 + 20 && x < X4 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y6 + 42 && y < Y6 + 48) :

             (array[235:232] == 4'b0110) ? (x > X4 + 20 && x < X4 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        
             (array[235:232] == 4'b0111) ?   (x > X4 + 20 && x < X4 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y6 + 12 && y < Y6 + 48) : 


             (array[235:232] == 4'b1000) ? (x > X4 + 20 && x < X4 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X4 + 45 && x < X4 + 52 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                         
             (array[235:232] == 4'b1001) ?  (x > X4 + 20 && x < X4 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                        (x > X4 + 20 && x < X4 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X4 + 45 && x < X4 + 52 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                        (x > X4 + 20 && x < X4 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        0;

assign num[59] = (array[239:236] == 4'b0001) ? (x > X5 + 30 && x < X5 + 42 && y > Y6 + 6 && y < Y6 + 48) :



              (array[239:236] == 4'b0010) ? ((x > X5 + 20 && x < X5 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y6 + 30 && y < Y6 + 42)) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y6 + 42 && y < Y6 + 48):


                
              (array[239:236] == 4'b0011) ? (x > X5 + 20 && x < X5 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y6 + 42 && y < Y6 + 48):

  
              (array[239:236] == 4'b0100) ? (x > X5 + 20 && x < X5 + 27 && y > Y6 + 6 && y < Y6 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y6 + 6 && y < Y6 + 48): 


             (array[239:236] == 4'b0101) ? (x > X5 + 20 && x < X5 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y6 + 42 && y < Y6 + 48) :

             (array[239:236] == 4'b0110) ? (x > X5 + 20 && x < X5 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        
             (array[239:236] == 4'b0111) ?   (x > X5 + 20 && x < X5 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y6 + 12 && y < Y6 + 48) : 


             (array[239:236] == 4'b1000) ? (x > X5 + 20 && x < X5 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X5 + 45 && x < X5 + 52 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                         
             (array[239:236] == 4'b1001) ?  (x > X5 + 20 && x < X5 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                        (x > X5 + 20 && x < X5 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X5 + 45 && x < X5 + 52 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                        (x > X5 + 20 && x < X5 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        0;

assign num[60] = (array[243:240] == 4'b0001) ? (x > X6 + 30 && x < X6 + 42 && y > Y6 + 6 && y < Y6 + 48) :



              (array[243:240] == 4'b0010) ? ((x > X6 + 20 && x < X6 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y6 + 30 && y < Y6 + 42)) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y6 + 42 && y < Y6 + 48):


                
              (array[243:240] == 4'b0011) ? (x > X6 + 20 && x < X6 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y6 + 42 && y < Y6 + 48):

  
              (array[243:240] == 4'b0100) ? (x > X6 + 20 && x < X6 + 27 && y > Y6 + 6 && y < Y6 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y6 + 6 && y < Y6 + 48): 


             (array[243:240] == 4'b0101) ? (x > X6 + 20 && x < X6 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y6 + 42 && y < Y6 + 48) :

             (array[243:240] == 4'b0110) ? (x > X6 + 20 && x < X6 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        
             (array[243:240] == 4'b0111) ?   (x > X6 + 20 && x < X6 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y6 + 12 && y < Y6 + 48) : 


             (array[243:240] == 4'b1000) ? (x > X6 + 20 && x < X6 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X6 + 45 && x < X6 + 52 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                         
             (array[243:240] == 4'b1001) ?  (x > X6 + 20 && x < X6 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                        (x > X6 + 20 && x < X6 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X6 + 45 && x < X6 + 52 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                        (x > X6 + 20 && x < X6 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        0;

assign num[61] = (array[247:244] == 4'b0001) ? (x > X7 + 30 && x < X7 + 42 && y > Y6 + 6 && y < Y6 + 48) :



              (array[247:244] == 4'b0010) ? ((x > X7 + 20 && x < X7 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y6 + 30 && y < Y6 + 42)) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y6 + 42 && y < Y6 + 48):


                
              (array[247:244] == 4'b0011) ? (x > X7 + 20 && x < X7 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y6 + 42 && y < Y6 + 48):

  
              (array[247:244] == 4'b0100) ? (x > X7 + 20 && x < X7 + 27 && y > Y6 + 6 && y < Y6 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y6 + 6 && y < Y6 + 48): 


             (array[247:244] == 4'b0101) ? (x > X7 + 20 && x < X7 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y6 + 42 && y < Y6 + 48) :

             (array[247:244] == 4'b0110) ? (x > X7 + 20 && x < X7 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        
             (array[247:244] == 4'b0111) ?   (x > X7 + 20 && x < X7 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y6 + 12 && y < Y6 + 48) : 


             (array[247:244] == 4'b1000) ? (x > X7 + 20 && x < X7 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X7 + 45 && x < X7 + 52 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                         
             (array[247:244] == 4'b1001) ?  (x > X7 + 20 && x < X7 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                        (x > X7 + 20 && x < X7 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X7 + 45 && x < X7 + 52 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                        (x > X7 + 20 && x < X7 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        0;

assign num[62] = (array[251:248] == 4'b0001) ? (x > X8 + 30 && x < X8 + 42 && y > Y6 + 6 && y < Y6 + 48) :



              (array[251:248] == 4'b0010) ? ((x > X8 + 20 && x < X8 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y6 + 30 && y < Y6 + 42)) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y6 + 42 && y < Y6 + 48):


                
              (array[251:248] == 4'b0011) ? (x > X8 + 20 && x < X8 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y6 + 12 && y < Y6 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y6 + 42 && y < Y6 + 48):

  
              (array[251:248] == 4'b0100) ? (x > X8 + 20 && x < X8 + 27 && y > Y6 + 6 && y < Y6 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y6 + 6 && y < Y6 + 48): 


             (array[251:248] == 4'b0101) ? (x > X8 + 20 && x < X8 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y6 + 42 && y < Y6 + 48) :

             (array[251:248] == 4'b0110) ? (x > X8 + 20 && x < X8 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y6 + 24 && y < Y6 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y6 + 30 && y < Y6 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        
             (array[251:248] == 4'b0111) ?   (x > X8 + 20 && x < X8 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y6 + 12 && y < Y6 + 48) : 


             (array[251:248] == 4'b1000) ? (x > X8 + 20 && x < X8 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X8 + 45 && x < X8 + 52 && y > Y6 + 12 && y < Y6 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                         
             (array[251:248] == 4'b1001) ?  (x > X8 + 20 && x < X8 + 52 && y > Y6 + 6 && y < Y6 + 12) || 
                                        (x > X8 + 20 && x < X8 + 27 && y > Y6 + 12 && y < Y6 + 24) || 
                                        (x > X8 + 45 && x < X8 + 52 && y > Y6 + 12 && y < Y6 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y6 + 24 && y < Y6 + 30) ||
                                        (x > X8 + 20 && x < X8 + 52 && y > Y6 + 42 && y < Y6 + 48) : 
                                        0;



assign num[63] = (array[255:252] == 4'b0001) ? (x > X0 + 30 && x < X0 + 42 && y > Y7 + 6 && y < Y7 + 48) :



              (array[255:252] == 4'b0010) ? ((x > X0 + 20 && x < X0 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y7 + 30 && y < Y7 + 42)) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y7 + 42 && y < Y7 + 48):


                
              (array[255:252] == 4'b0011) ? (x > X0 + 20 && x < X0 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y7 + 42 && y < Y7 + 48):

  
              (array[255:252] == 4'b0100) ? (x > X0 + 20 && x < X0 + 27 && y > Y7 + 6 && y < Y7 + 24) || 
                                       (x > X0 + 20 && x < X0 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X0 + 45 && x < X0 + 52 && y > Y7 + 6 && y < Y7 + 48): 


             (array[255:252] == 4'b0101) ? (x > X0 + 20 && x < X0 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y7 + 42 && y < Y7 + 48) :

             (array[255:252] == 4'b0110) ? (x > X0 + 20 && x < X0 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X0 + 20 && x < X0 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        
             (array[255:252] == 4'b0111) ?   (x > X0 + 20 && x < X0 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                         (x > X0 + 45 && x < X0 + 52 && y > Y7 + 12 && y < Y7 + 48) : 


             (array[255:252] == 4'b1000) ? (x > X0 + 20 && x < X0 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X0 + 20 && x < X0 + 27 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X0 + 45 && x < X0 + 52 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                       (x > X0 + 20 && x < X0 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                         
             (array[255:252] == 4'b1001) ?  (x > X0 + 20 && x < X0 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                        (x > X0 + 20 && x < X0 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X0 + 45 && x < X0 + 52 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X0 + 20 && x < X0 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                        (x > X0 + 20 && x < X0 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        0;

assign num[64] = (array[259:256] == 4'b0001) ? (x > X1 + 30 && x < X1 + 42 && y > Y7 + 6 && y < Y7 + 48) :



              (array[259:256] == 4'b0010) ? ((x > X1 + 20 && x < X1 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y7 + 30 && y < Y7 + 42)) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y7 + 42 && y < Y7 + 48):


                
              (array[259:256] == 4'b0011) ? (x > X1 + 20 && x < X1 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y7 + 42 && y < Y7 + 48):

  
              (array[259:256] == 4'b0100) ? (x > X1 + 20 && x < X1 + 27 && y > Y7 + 6 && y < Y7 + 24) || 
                                       (x > X1 + 20 && x < X1 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X1 + 45 && x < X1 + 52 && y > Y7 + 6 && y < Y7 + 48): 


             (array[259:256] == 4'b0101) ? (x > X1 + 20 && x < X1 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y7 + 42 && y < Y7 + 48) :

             (array[259:256] == 4'b0110) ? (x > X1 + 20 && x < X1 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X1 + 20 && x < X1 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        
             (array[259:256] == 4'b0111) ?   (x > X1 + 20 && x < X1 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                         (x > X1 + 45 && x < X1 + 52 && y > Y7 + 12 && y < Y7 + 48) : 


             (array[259:256] == 4'b1000) ? (x > X1 + 20 && x < X1 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X1 + 20 && x < X1 + 27 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X1 + 45 && x < X1 + 52 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                       (x > X1 + 20 && x < X1 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                         
             (array[259:256] == 4'b1001) ?  (x > X1 + 20 && x < X1 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                        (x > X1 + 20 && x < X1 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X1 + 45 && x < X1 + 52 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X1 + 20 && x < X1 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                        (x > X1 + 20 && x < X1 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        0;

assign num[65] = (array[263:260] == 4'b0001) ? (x > X2 + 30 && x < X2 + 42 && y > Y7 + 6 && y < Y7 + 48) :



              (array[263:260] == 4'b0010) ? ((x > X2 + 20 && x < X2 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y7 + 30 && y < Y7 + 42)) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y7 + 42 && y < Y7 + 48):


                
              (array[263:260] == 4'b0011) ? (x > X2 + 20 && x < X2 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y7 + 42 && y < Y7 + 48):

  
              (array[263:260] == 4'b0100) ? (x > X2 + 20 && x < X2 + 27 && y > Y7 + 6 && y < Y7 + 24) || 
                                       (x > X2 + 20 && x < X2 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X2 + 45 && x < X2 + 52 && y > Y7 + 6 && y < Y7 + 48): 


             (array[263:260] == 4'b0101) ? (x > X2 + 20 && x < X2 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y7 + 42 && y < Y7 + 48) :

             (array[263:260] == 4'b0110) ? (x > X2 + 20 && x < X2 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X2 + 20 && x < X2 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        
             (array[263:260] == 4'b0111) ?   (x > X2 + 20 && x < X2 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                         (x > X2 + 45 && x < X2 + 52 && y > Y7 + 12 && y < Y7 + 48) : 


             (array[263:260] == 4'b1000) ? (x > X2 + 20 && x < X2 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X2 + 20 && x < X2 + 27 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X2 + 45 && x < X2 + 52 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                       (x > X2 + 20 && x < X2 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                         
             (array[263:260] == 4'b1001) ?  (x > X2 + 20 && x < X2 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                        (x > X2 + 20 && x < X2 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X2 + 45 && x < X2 + 52 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X2 + 20 && x < X2 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                        (x > X2 + 20 && x < X2 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        0;


assign num[66] = (array[267:264] == 4'b0001) ? (x > X3 + 30 && x < X3 + 42 && y > Y7 + 6 && y < Y7 + 48) :



              (array[267:264] == 4'b0010) ? ((x > X3 + 20 && x < X3 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y7 + 30 && y < Y7 + 42)) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y7 + 42 && y < Y7 + 48):


                
              (array[267:264] == 4'b0011) ? (x > X3 + 20 && x < X3 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y7 + 42 && y < Y7 + 48):

  
              (array[267:264] == 4'b0100) ? (x > X3 + 20 && x < X3 + 27 && y > Y7 + 6 && y < Y7 + 24) || 
                                       (x > X3 + 20 && x < X3 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X3 + 45 && x < X3 + 52 && y > Y7 + 6 && y < Y7 + 48): 


             (array[267:264] == 4'b0101) ? (x > X3 + 20 && x < X3 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y7 + 42 && y < Y7 + 48) :

             (array[267:264] == 4'b0110) ? (x > X3 + 20 && x < X3 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X3 + 20 && x < X3 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        
             (array[267:264] == 4'b0111) ?   (x > X3 + 20 && x < X3 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                         (x > X3 + 45 && x < X3 + 52 && y > Y7 + 12 && y < Y7 + 48) : 


             (array[267:264] == 4'b1000) ? (x > X3 + 20 && x < X3 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X3 + 20 && x < X3 + 27 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X3 + 45 && x < X3 + 52 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                       (x > X3 + 20 && x < X3 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                         
             (array[267:264] == 4'b1001) ?  (x > X3 + 20 && x < X3 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                        (x > X3 + 20 && x < X3 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X3 + 45 && x < X3 + 52 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X3 + 20 && x < X3 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                        (x > X3 + 20 && x < X3 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        0;


assign num[67] = (array[271:268] == 4'b0001) ? (x > X4 + 30 && x < X4 + 42 && y > Y7 + 6 && y < Y7 + 48) :



              (array[271:268] == 4'b0010) ? ((x > X4 + 20 && x < X4 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y7 + 30 && y < Y7 + 42)) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y7 + 42 && y < Y7 + 48):


                
              (array[271:268] == 4'b0011) ? (x > X4 + 20 && x < X4 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y7 + 42 && y < Y7 + 48):

  
              (array[271:268] == 4'b0100) ? (x > X4 + 20 && x < X4 + 27 && y > Y7 + 6 && y < Y7 + 24) || 
                                       (x > X4 + 20 && x < X4 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X4 + 45 && x < X4 + 52 && y > Y7 + 6 && y < Y7 + 48): 


             (array[271:268] == 4'b0101) ? (x > X4 + 20 && x < X4 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y7 + 42 && y < Y7 + 48) :

             (array[271:268] == 4'b0110) ? (x > X4 + 20 && x < X4 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X4 + 20 && x < X4 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        
             (array[271:268] == 4'b0111) ?   (x > X4 + 20 && x < X4 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                         (x > X4 + 45 && x < X4 + 52 && y > Y7 + 12 && y < Y7 + 48) : 


             (array[271:268] == 4'b1000) ? (x > X4 + 20 && x < X4 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X4 + 20 && x < X4 + 27 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X4 + 45 && x < X4 + 52 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                       (x > X4 + 20 && x < X4 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                         
             (array[271:268] == 4'b1001) ?  (x > X4 + 20 && x < X4 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                        (x > X4 + 20 && x < X4 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X4 + 45 && x < X4 + 52 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X4 + 20 && x < X4 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                        (x > X4 + 20 && x < X4 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        0;

assign num[68] = (array[275:272] == 4'b0001) ? (x > X5 + 30 && x < X5 + 42 && y > Y7 + 6 && y < Y7 + 48) :



              (array[275:272] == 4'b0010) ? ((x > X5 + 20 && x < X5 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y7 + 30 && y < Y7 + 42)) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y7 + 42 && y < Y7 + 48):


                
              (array[275:272] == 4'b0011) ? (x > X5 + 20 && x < X5 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y7 + 42 && y < Y7 + 48):

  
              (array[275:272] == 4'b0100) ? (x > X5 + 20 && x < X5 + 27 && y > Y7 + 6 && y < Y7 + 24) || 
                                       (x > X5 + 20 && x < X5 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X5 + 45 && x < X5 + 52 && y > Y7 + 6 && y < Y7 + 48): 


             (array[275:272] == 4'b0101) ? (x > X5 + 20 && x < X5 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y7 + 42 && y < Y7 + 48) :

             (array[275:272] == 4'b0110) ? (x > X5 + 20 && x < X5 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X5 + 20 && x < X5 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        
             (array[275:272] == 4'b0111) ?   (x > X5 + 20 && x < X5 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                         (x > X5 + 45 && x < X5 + 52 && y > Y7 + 12 && y < Y7 + 48) : 


             (array[275:272] == 4'b1000) ? (x > X5 + 20 && x < X5 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X5 + 20 && x < X5 + 27 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X5 + 45 && x < X5 + 52 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                       (x > X5 + 20 && x < X5 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                         
             (array[275:272] == 4'b1001) ?  (x > X5 + 20 && x < X5 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                        (x > X5 + 20 && x < X5 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X5 + 45 && x < X5 + 52 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X5 + 20 && x < X5 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                        (x > X5 + 20 && x < X5 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        0;

assign num[69] = (array[279:276] == 4'b0001) ? (x > X6 + 30 && x < X6 + 42 && y > Y7 + 6 && y < Y7 + 48) :



              (array[279:276] == 4'b0010) ? ((x > X6 + 20 && x < X6 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y7 + 30 && y < Y7 + 42)) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y7 + 42 && y < Y7 + 48):


                
              (array[279:276] == 4'b0011) ? (x > X6 + 20 && x < X6 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y7 + 42 && y < Y7 + 48):

  
              (array[279:276] == 4'b0100) ? (x > X6 + 20 && x < X6 + 27 && y > Y7 + 6 && y < Y7 + 24) || 
                                       (x > X6 + 20 && x < X6 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X6 + 45 && x < X6 + 52 && y > Y7 + 6 && y < Y7 + 48): 


             (array[279:276] == 4'b0101) ? (x > X6 + 20 && x < X6 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y7 + 42 && y < Y7 + 48) :

             (array[279:276] == 4'b0110) ? (x > X6 + 20 && x < X6 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X6 + 20 && x < X6 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        
             (array[279:276] == 4'b0111) ?   (x > X6 + 20 && x < X6 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                         (x > X6 + 45 && x < X6 + 52 && y > Y7 + 12 && y < Y7 + 48) : 


             (array[279:276] == 4'b1000) ? (x > X6 + 20 && x < X6 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X6 + 20 && x < X6 + 27 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X6 + 45 && x < X6 + 52 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                       (x > X6 + 20 && x < X6 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                         
             (array[279:276] == 4'b1001) ?  (x > X6 + 20 && x < X6 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                        (x > X6 + 20 && x < X6 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X6 + 45 && x < X6 + 52 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X6 + 20 && x < X6 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                        (x > X6 + 20 && x < X6 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        0;

assign num[70] = (array[283:280] == 4'b0001) ? (x > X7 + 30 && x < X7 + 42 && y > Y7 + 6 && y < Y7 + 48) :



              (array[283:280] == 4'b0010) ? ((x > X7 + 20 && x < X7 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y7 + 30 && y < Y7 + 42)) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y7 + 42 && y < Y7 + 48):


                
              (array[283:280] == 4'b0011) ? (x > X7 + 20 && x < X7 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y7 + 42 && y < Y7 + 48):

  
              (array[283:280] == 4'b0100) ? (x > X7 + 20 && x < X7 + 27 && y > Y7 + 6 && y < Y7 + 24) || 
                                       (x > X7 + 20 && x < X7 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X7 + 45 && x < X7 + 52 && y > Y7 + 6 && y < Y7 + 48): 


             (array[283:280] == 4'b0101) ? (x > X7 + 20 && x < X7 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y7 + 42 && y < Y7 + 48) :

             (array[283:280] == 4'b0110) ? (x > X7 + 20 && x < X7 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X7 + 20 && x < X7 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        
             (array[283:280] == 4'b0111) ?   (x > X7 + 20 && x < X7 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                         (x > X7 + 45 && x < X7 + 52 && y > Y7 + 12 && y < Y7 + 48) : 


             (array[283:280] == 4'b1000) ? (x > X7 + 20 && x < X7 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X7 + 20 && x < X7 + 27 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X7 + 45 && x < X7 + 52 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                       (x > X7 + 20 && x < X7 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                         
             (array[283:280] == 4'b1001) ?  (x > X7 + 20 && x < X7 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                        (x > X7 + 20 && x < X7 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X7 + 45 && x < X7 + 52 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X7 + 20 && x < X7 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                        (x > X7 + 20 && x < X7 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        0;

assign num[71] = (array[287:284] == 4'b0001) ? (x > X8 + 30 && x < X8 + 42 && y > Y7 + 6 && y < Y7 + 48) :



              (array[287:284] == 4'b0010) ? ((x > X8 + 20 && x < X8 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y7 + 30 && y < Y7 + 42)) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y7 + 42 && y < Y7 + 48):


                
              (array[287:284] == 4'b0011) ? (x > X8 + 20 && x < X8 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y7 + 12 && y < Y7 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y7 + 42 && y < Y7 + 48):

  
              (array[287:284] == 4'b0100) ? (x > X8 + 20 && x < X8 + 27 && y > Y7 + 6 && y < Y7 + 24) || 
                                       (x > X8 + 20 && x < X8 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                       (x > X8 + 45 && x < X8 + 52 && y > Y7 + 6 && y < Y7 + 48): 


             (array[287:284] == 4'b0101) ? (x > X8 + 20 && x < X8 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y7 + 42 && y < Y7 + 48) :

             (array[287:284] == 4'b0110) ? (x > X8 + 20 && x < X8 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y7 + 24 && y < Y7 + 30) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y7 + 30 && y < Y7 + 42) ||
                                         (x > X8 + 20 && x < X8 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        
             (array[287:284] == 4'b0111) ?   (x > X8 + 20 && x < X8 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                         (x > X8 + 45 && x < X8 + 52 && y > Y7 + 12 && y < Y7 + 48) : 


             (array[287:284] == 4'b1000) ? (x > X8 + 20 && x < X8 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                       (x > X8 + 20 && x < X8 + 27 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X8 + 45 && x < X8 + 52 && y > Y7 + 12 && y < Y7 + 42) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                       (x > X8 + 20 && x < X8 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                         
             (array[287:284] == 4'b1001) ?  (x > X8 + 20 && x < X8 + 52 && y > Y7 + 6 && y < Y7 + 12) || 
                                        (x > X8 + 20 && x < X8 + 27 && y > Y7 + 12 && y < Y7 + 24) || 
                                        (x > X8 + 45 && x < X8 + 52 && y > Y7 + 12 && y < Y7 + 42) || 
                                        (x > X8 + 20 && x < X8 + 52 && y > Y7 + 24 && y < Y7 + 30) ||
                                        (x > X8 + 20 && x < X8 + 52 && y > Y7 + 42 && y < Y7 + 48) : 
                                        0;
                                        

      
                
  
  
                
                
                
                
                
endmodule
